//fn6

	`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   12:10:21 10/01/2015
// Design Name:   prof_test
// Module Name:   D:/Pavan_FPGA_Projects/cam_test_1/tb.v
// Project Name:  cam_test_1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: prof_test
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb;

	// Inputs
	reg clk;
	reg reset;
	reg [0:31] P_Trace_Instruction;
	reg [0:31] P_Trace_PC;
	reg P_Trace_Valid_Instr;
	reg P_Trace_Jump_Taken;
	
	reg sel;
	reg [4:0] in_addr;

	// Outputs
	//wire [3:0] match_addr;
	//wire busy;
	//wire [31:0] P_Count;
	wire [31:0] data_out;
   //wire [31:0] final_cnt;
	// Instantiate the Unit Under Test (UUT)
	f_l_prof uut (
		.clk(clk), 
		.reset(reset), 
		.P_Trace_Instruction(P_Trace_Instruction), 
		.P_Trace_PC(P_Trace_PC), 
		.P_Trace_Valid_Instr(P_Trace_Valid_Instr), 
		.P_Trace_Jump_Taken(P_Trace_Jump_Taken)
		//.match_addr(match_addr),
		//.busy(busy),
		//.sel(sel),
		//.in_addr(in_addr),
		//.data_out(data_out)
		//.final_cnt(final_cnt)
	);




initial
begin
/*$monitor ("time=%d,pc=%h,loop_det=%b,jmp_taken=%b, match= %b, temp_pc= %h ,state =%b, cnt_enable = %b, we = %b ,load =%b,clear =%b,busy =%b, count =%h,addr =%b, match_addr=%b, write_en= %b , data_out = %h, mux_addr = %b, sel=%b, ram_data_in= %h",
$time,P_Trace_PC,uut.loop_det,P_Trace_Jump_Taken,uut.cam_match,uut.temp_pc,uut.state,uut.cnt_enable,uut.cam_we,uut.load,uut.clear,uut.cam_busy,uut.P_Count,uut.addr,uut.match_addr,uut.write_en,uut.data_out,uut.mux_addr,uut.sel,uut.ram_data_in);
*/
/*M
$monitor ("time=%d,pc=%h,P_Trace_Valid_Instr=%b, P_Trace_Instruction=%h, loop_det=%b,jmp_taken=%b, match= %b, temp_pc= %h ,state =%d,count =%h,addr =%b, match_addr=%b, write_en= %b , data_out = %h, mux_addr = %b,ram_data_in= %h",
$time,P_Trace_PC,P_Trace_Valid_Instr,P_Trace_Instruction, uut.loop_det,P_Trace_Jump_Taken,uut.cam_match,uut.temp_pc,uut.state,uut.P_Count,uut.addr,uut.match_addr,uut.write_en,uut.data_out,uut.mux_addr,uut.ram_data_in);
*/
/*
$monitor ("time=%d,pc=%h,P_Trace_Valid_Instr=%b, P_Trace_Instruction=%h, cam_busy=%b, cam_we=%b, loop_det=%b,jmp_taken=%b, match= %b, load=%b, cnt_enable=%b, addr_cnt_enable=%b, temp_pc= %h ,state =%d, next_state =%d,count =%h,addr =%b, match_addr=%b, write_en= %b , data_out = %h, mux_addr = %b,ram_data_in= %h",
$time,P_Trace_PC,P_Trace_Valid_Instr,P_Trace_Instruction, uut.cam_busy, uut.cam_we, uut.loop_det,P_Trace_Jump_Taken,uut.cam_match,uut.load, uut.cnt_enable, uut.addr_cnt_enable,uut.temp_pc,uut.state,uut.next_state, uut.P_Count,uut.addr,uut.match_addr,uut.write_en,uut.data_out,uut.mux_addr,uut.ram_data_in);

*/
/*
$monitor ("t=%d,pc=%h,Valid_Instr=%b,P_Trace_Instr=%h, loop_det=%b,jmp_taken=%b, cnt_en=%b,ps=%d,ns=%d, p_count =%h, cam_busy=%b, cam_we=%b, match1=%b, match= %b, load=%b,  addr_cnt_enable=%b, temp_pc= %h ,addr =%b, cam_en= %b, match_addr=%b, sel_match=%b, cam_addr=%b, cam_addr_previous=%b, write_en= %b , data_out = %h, mux_addr = %b,ram_data_in= %h, f_Valid_Instr=%b, f_P_Trace_Jump_Taken=%b, f_loop_det=%b, i2=%b, flag_reg=%b, match_addr_RAM=%b, match_previous_addr=%b, final_cnt=%b flag_en=%b",
$time,P_Trace_PC,P_Trace_Valid_Instr,P_Trace_Instruction,uut.loop_det,P_Trace_Jump_Taken,uut.cnt_enable,uut.state,uut.next_state,uut.P_Count,uut.cam_busy,uut.cam_we,uut.cam_match1,uut.cam_match,uut.load,uut.addr_cnt_enable,uut.temp_pc,uut.addr, uut.cam_en, uut.match_addr, uut.sel_match, uut.cam_addr, uut.cam_addr_previous, uut.write_en,uut.data_out,uut.mux_addr,uut.ram_data_in, uut.f_Valid_Instr, uut.f_P_Trace_Jump_Taken, uut.f_loop_det, uut.i2, uut.flag_reg, uut.match_addr_RAM, uut.match_previous_addr, uut.final_cnt, uut.flag_en);
*/
/*$monitor ("t=%d,pc=%h,Valid_Instr=%b,P_Trace_Instr=%h, loop_det=%b,jmp_taken=%b, cnt_en=%b,ps=%d,ns=%d, p_count =%h, cam_we=%b,  match= %b, load=%b,  addr_cnt_enable=%b, temp_pc= %h ,addr =%b, cam_en= %b, match_addr=%b, write_en= %b , data_out = %h, mux_addr = %b,ram_data_in= %h, f_Valid_Instr=%b, f_P_Trace_Jump_Taken=%b, f_loop_det=%b, i2=%b, flag_reg=%b, match_addr_RAM=%b, match_previous_addr=%b, final_cnt=%b flag_en=%b",
$time,P_Trace_PC,P_Trace_Valid_Instr,P_Trace_Instruction,uut.loop_det,P_Trace_Jump_Taken,uut.cnt_enable,uut.state,uut.next_state,uut.P_Count,uut.cam_we,uut.cam_match,uut.load,uut.addr_cnt_enable,uut.temp_pc,uut.addr, uut.cam_en, uut.match_addr, uut.write_en,uut.data_out,uut.mux_addr,uut.ram_data_in, uut.f_Valid_Instr, uut.f_P_Trace_Jump_Taken, uut.f_loop_det, uut.i2, uut.flag_reg, uut.match_addr_RAM, uut.match_previous_addr, uut.final_cnt, uut.flag_en);

*/
sel = 1'b0;
in_addr = 4'b0000;

// will have to initialise//


#0 P_Trace_PC = 32'h00000124;
reset = 1'b0;
P_Trace_Instruction = 32'hFA61000C;
P_Trace_Valid_Instr = 1'b1;
clk = 1'b1;
sel = 1'b0;
in_addr = 4'b0000;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000184;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F40158;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000188;
reset = 1'b0;
P_Trace_Instruction = 32'h20A00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000188;
reset = 1'b0;
P_Trace_Instruction = 32'h20A00000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002DC;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFE0;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002E4;
reset = 1'b0;
P_Trace_Instruction = 32'hFA61001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002E8;
reset = 1'b0;
P_Trace_Instruction = 32'h12610000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002F0;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002F4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002F8;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F4FF94;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000002FC;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002FC;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000028C;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFE0;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000290;
reset = 1'b0;
P_Trace_Instruction = 32'hF9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000294;
reset = 1'b0;
P_Trace_Instruction = 32'hFA61001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000298;
reset = 1'b0;
P_Trace_Instruction = 32'h12610000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000029C;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F4FF14;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000002A0;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002A0;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001B0;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFF4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001B4;
reset = 1'b0;
P_Trace_Instruction = 32'hFA610008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001B8;
reset = 1'b0;
P_Trace_Instruction = 32'h12610000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001BC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8130004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C0;
reset = 1'b0;
P_Trace_Instruction = 32'hB800001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E4;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E8;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E4;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E8;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E4;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E8;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E4;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E8;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E4;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E8;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001C8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E0;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E4;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001E8;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001F0;
reset = 1'b0;
P_Trace_Instruction = 32'h10330000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001F4;
reset = 1'b0;
P_Trace_Instruction = 32'hEA610008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001F8;
reset = 1'b0;
P_Trace_Instruction = 32'h3021000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001FC;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000200;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000200;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002A4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8600814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002A8;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F4FF5C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000002AC;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002AC;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000204;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFF4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000208;
reset = 1'b0;
P_Trace_Instruction = 32'hFA610008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000020C;
reset = 1'b0;
P_Trace_Instruction = 32'h12610000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000210;
reset = 1'b0;
P_Trace_Instruction = 32'hF8130004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000214;
reset = 1'b0;
P_Trace_Instruction = 32'hB800001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000230;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000238;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000023C;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000021C;
reset = 1'b0;
P_Trace_Instruction = 32'h3063FFFF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000220;
reset = 1'b0;
P_Trace_Instruction = 32'hF86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000228;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000022C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000230;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000238;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000023C;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000021C;
reset = 1'b0;
P_Trace_Instruction = 32'h3063FFFF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000220;
reset = 1'b0;
P_Trace_Instruction = 32'hF86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000228;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000022C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000230;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000238;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000023C;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000021C;
reset = 1'b0;
P_Trace_Instruction = 32'h3063FFFF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000220;
reset = 1'b0;
P_Trace_Instruction = 32'hF86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000228;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000022C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000230;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000238;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000023C;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000021C;
reset = 1'b0;
P_Trace_Instruction = 32'h3063FFFF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000220;
reset = 1'b0;
P_Trace_Instruction = 32'hF86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000228;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000022C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000230;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000238;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000023C;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000218;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000021C;
reset = 1'b0;
P_Trace_Instruction = 32'h3063FFFF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000220;
reset = 1'b0;
P_Trace_Instruction = 32'hF86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000224;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000228;
reset = 1'b0;
P_Trace_Instruction = 32'h30630001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000022C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000230;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000234;
reset = 1'b0;
P_Trace_Instruction = 32'h32400004;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000238;
reset = 1'b0;
P_Trace_Instruction = 32'h16439001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000023C;
reset = 1'b0;
P_Trace_Instruction = 32'hBCB2FFDC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000240;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000244;
reset = 1'b0;
P_Trace_Instruction = 32'h10330000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000248;
reset = 1'b0;
P_Trace_Instruction = 32'hEA610008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000024C;
reset = 1'b0;
P_Trace_Instruction = 32'h3021000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000250;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000254;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000254;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002B0;
reset = 1'b0;
P_Trace_Instruction = 32'hF86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002B4;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F4FFA4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000002B8;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002B8;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000258;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFF4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000025C;
reset = 1'b0;
P_Trace_Instruction = 32'hFA610008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000260;
reset = 1'b0;
P_Trace_Instruction = 32'h12610000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000264;
reset = 1'b0;
P_Trace_Instruction = 32'hE8800814;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000268;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000268;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000268;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000026C;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000270;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000274;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000278;
reset = 1'b0;
P_Trace_Instruction = 32'h10330000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000027C;
reset = 1'b0;
P_Trace_Instruction = 32'hEA610008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000280;
reset = 1'b0;
P_Trace_Instruction = 32'h3021000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000284;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000288;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000288;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002BC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8600818;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8600818;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10330000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002CC;
reset = 1'b0;
P_Trace_Instruction = 32'hEA61001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002D0;
reset = 1'b0;
P_Trace_Instruction = 32'h30210020;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002D4;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000002D8;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000002D8;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000300;
reset = 1'b0;
P_Trace_Instruction = 32'hF8600818;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000304;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000308;
reset = 1'b0;
P_Trace_Instruction = 32'hE9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000030C;
reset = 1'b0;
P_Trace_Instruction = 32'h10330000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000310;
reset = 1'b0;
P_Trace_Instruction = 32'hEA61001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000314;
reset = 1'b0;
P_Trace_Instruction = 32'h30210020;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000318;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h0000031C;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000031C;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000018C;
reset = 1'b0;
P_Trace_Instruction = 32'h32630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000190;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F40510;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000194;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000194;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000006A0;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFF8;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000006A4;
reset = 1'b0;
P_Trace_Instruction = 32'hD9E00800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000006A8;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F4F9C8;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000006AC;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000006AC;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000070;
reset = 1'b0;
P_Trace_Instruction = 32'hE06007F8;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000074;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFE4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000074;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFE4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000078;
reset = 1'b0;
P_Trace_Instruction = 32'hBE03001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h0000007C;
reset = 1'b0;
P_Trace_Instruction = 32'hF9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000007C;
reset = 1'b0;
P_Trace_Instruction = 32'hF9E10000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000094;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D0;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000094;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D0;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000094;
reset = 1'b0;
P_Trace_Instruction = 32'hE86006D0;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000098;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000098;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000098;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000009C;
reset = 1'b0;
P_Trace_Instruction = 32'hBE24FFEC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000A0;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000A4;
reset = 1'b0;
P_Trace_Instruction = 32'hB0000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000A8;
reset = 1'b0;
P_Trace_Instruction = 32'h30600000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000AC;
reset = 1'b0;
P_Trace_Instruction = 32'hBC030010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000000B0;
reset = 1'b0;
P_Trace_Instruction = 32'h30A007EC;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000B0;
reset = 1'b0;
P_Trace_Instruction = 32'h30A007EC;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000BC;
reset = 1'b0;
P_Trace_Instruction = 32'h30600001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C0;
reset = 1'b0;
P_Trace_Instruction = 32'hF06007F8;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE9E10000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE9E10000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C8;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000000CC;
reset = 1'b0;
P_Trace_Instruction = 32'h3021001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000CC;
reset = 1'b0;
P_Trace_Instruction = 32'h3021001C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000006B0;
reset = 1'b0;
P_Trace_Instruction = 32'hC9E00800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000006B0;
reset = 1'b0;
P_Trace_Instruction = 32'hC9E00800;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000006B0;
reset = 1'b0;
P_Trace_Instruction = 32'hC9E00800;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000006B4;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000006B8;
reset = 1'b0;
P_Trace_Instruction = 32'h30210008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000006B8;
reset = 1'b0;
P_Trace_Instruction = 32'h30210008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000198;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F40190;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h0000019C;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000019C;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000328;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h0000032C;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000032C;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001A0;
reset = 1'b0;
P_Trace_Instruction = 32'hC9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001A4;
reset = 1'b0;
P_Trace_Instruction = 32'h30730000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001A4;
reset = 1'b0;
P_Trace_Instruction = 32'h30730000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001A8;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000001AC;
reset = 1'b0;
P_Trace_Instruction = 32'h20210014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001AC;
reset = 1'b0;
P_Trace_Instruction = 32'h20210014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000064;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F403BC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000068;
reset = 1'b0;
P_Trace_Instruction = 32'h30A30000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000068;
reset = 1'b0;
P_Trace_Instruction = 32'h30A30000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000420;
reset = 1'b0;
P_Trace_Instruction = 32'hBA0C0018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;



//$display("ram_out=%h",uut.ram_out);
    $finish;
end

always
#10 clk=~clk;



	
      
endmodule