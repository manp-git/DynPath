//bcnt

	`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   12:10:21 10/01/2015
// Design Name:   prof_test
// Module Name:   D:/Pavan_FPGA_Projects/cam_test_1/tb.v
// Project Name:  cam_test_1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: prof_test
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb;

	// Inputs
	reg clk;
	reg reset;
	reg [0:31] P_Trace_Instruction;
	reg [0:31] P_Trace_PC;
	reg P_Trace_Valid_Instr;
	reg P_Trace_Jump_Taken;
	
	reg sel;
	reg [4:0] in_addr;

	// Outputs
	//wire [3:0] match_addr;
	//wire busy;
	//wire [31:0] P_Count;
	wire [31:0] data_out;
   //wire [31:0] final_cnt;
	// Instantiate the Unit Under Test (UUT)
	f_l_prof uut (
		.clk(clk), 
		.reset(reset), 
		.P_Trace_Instruction(P_Trace_Instruction), 
		.P_Trace_PC(P_Trace_PC), 
		.P_Trace_Valid_Instr(P_Trace_Valid_Instr), 
		.P_Trace_Jump_Taken(P_Trace_Jump_Taken)
		//.match_addr(match_addr),
		//.busy(busy),
		//.sel(sel),
		//.in_addr(in_addr),
		//.data_out(data_out)
		//.final_cnt(final_cnt)
	);




initial
begin
/*$monitor ("time=%d,pc=%h,loop_det=%b,jmp_taken=%b, match= %b, temp_pc= %h ,state =%b, cnt_enable = %b, we = %b ,load =%b,clear =%b,busy =%b, count =%h,addr =%b, match_addr=%b, write_en= %b , data_out = %h, mux_addr = %b, sel=%b, ram_data_in= %h",
$time,P_Trace_PC,uut.loop_det,P_Trace_Jump_Taken,uut.cam_match,uut.temp_pc,uut.state,uut.cnt_enable,uut.cam_we,uut.load,uut.clear,uut.cam_busy,uut.P_Count,uut.addr,uut.match_addr,uut.write_en,uut.data_out,uut.mux_addr,uut.sel,uut.ram_data_in);
*/
/*M
$monitor ("time=%d,pc=%h,P_Trace_Valid_Instr=%b, P_Trace_Instruction=%h, loop_det=%b,jmp_taken=%b, match= %b, temp_pc= %h ,state =%d,count =%h,addr =%b, match_addr=%b, write_en= %b , data_out = %h, mux_addr = %b,ram_data_in= %h",
$time,P_Trace_PC,P_Trace_Valid_Instr,P_Trace_Instruction, uut.loop_det,P_Trace_Jump_Taken,uut.cam_match,uut.temp_pc,uut.state,uut.P_Count,uut.addr,uut.match_addr,uut.write_en,uut.data_out,uut.mux_addr,uut.ram_data_in);
*/
/*
$monitor ("time=%d,pc=%h,P_Trace_Valid_Instr=%b, P_Trace_Instruction=%h, cam_busy=%b, cam_we=%b, loop_det=%b,jmp_taken=%b, match= %b, load=%b, cnt_enable=%b, addr_cnt_enable=%b, temp_pc= %h ,state =%d, next_state =%d,count =%h,addr =%b, match_addr=%b, write_en= %b , data_out = %h, mux_addr = %b,ram_data_in= %h",
$time,P_Trace_PC,P_Trace_Valid_Instr,P_Trace_Instruction, uut.cam_busy, uut.cam_we, uut.loop_det,P_Trace_Jump_Taken,uut.cam_match,uut.load, uut.cnt_enable, uut.addr_cnt_enable,uut.temp_pc,uut.state,uut.next_state, uut.P_Count,uut.addr,uut.match_addr,uut.write_en,uut.data_out,uut.mux_addr,uut.ram_data_in);

*/
/*
$monitor ("t=%d,pc=%h,Valid_Instr=%b,P_Trace_Instr=%h, loop_det=%b,jmp_taken=%b, cnt_en=%b,ps=%d,ns=%d, p_count =%h, cam_busy=%b, cam_we=%b, match1=%b, match= %b, load=%b,  addr_cnt_enable=%b, temp_pc= %h ,addr =%b, cam_en= %b, match_addr=%b, sel_match=%b, cam_addr=%b, cam_addr_previous=%b, write_en= %b , data_out = %h, mux_addr = %b,ram_data_in= %h, f_Valid_Instr=%b, f_P_Trace_Jump_Taken=%b, f_loop_det=%b, i2=%b, flag_reg=%b, match_addr_RAM=%b, match_previous_addr=%b, final_cnt=%b flag_en=%b",
$time,P_Trace_PC,P_Trace_Valid_Instr,P_Trace_Instruction,uut.loop_det,P_Trace_Jump_Taken,uut.cnt_enable,uut.state,uut.next_state,uut.P_Count,uut.cam_busy,uut.cam_we,uut.cam_match1,uut.cam_match,uut.load,uut.addr_cnt_enable,uut.temp_pc,uut.addr, uut.cam_en, uut.match_addr, uut.sel_match, uut.cam_addr, uut.cam_addr_previous, uut.write_en,uut.data_out,uut.mux_addr,uut.ram_data_in, uut.f_Valid_Instr, uut.f_P_Trace_Jump_Taken, uut.f_loop_det, uut.i2, uut.flag_reg, uut.match_addr_RAM, uut.match_previous_addr, uut.final_cnt, uut.flag_en);
*/
/*$monitor ("t=%d,pc=%h,Valid_Instr=%b,P_Trace_Instr=%h, loop_det=%b,jmp_taken=%b, cnt_en=%b,ps=%d,ns=%d, p_count =%h, cam_we=%b,  match= %b, load=%b,  addr_cnt_enable=%b, temp_pc= %h ,addr =%b, cam_en= %b, match_addr=%b, write_en= %b , data_out = %h, mux_addr = %b,ram_data_in= %h, f_Valid_Instr=%b, f_P_Trace_Jump_Taken=%b, f_loop_det=%b, i2=%b, flag_reg=%b, match_addr_RAM=%b, match_previous_addr=%b, final_cnt=%b flag_en=%b",
$time,P_Trace_PC,P_Trace_Valid_Instr,P_Trace_Instruction,uut.loop_det,P_Trace_Jump_Taken,uut.cnt_enable,uut.state,uut.next_state,uut.P_Count,uut.cam_we,uut.cam_match,uut.load,uut.addr_cnt_enable,uut.temp_pc,uut.addr, uut.cam_en, uut.match_addr, uut.write_en,uut.data_out,uut.mux_addr,uut.ram_data_in, uut.f_Valid_Instr, uut.f_P_Trace_Jump_Taken, uut.f_loop_det, uut.i2, uut.flag_reg, uut.match_addr_RAM, uut.match_previous_addr, uut.final_cnt, uut.flag_en);

*/
sel = 1'b0;
in_addr = 4'b0000;

// will have to initialise//


#0 P_Trace_PC = 32'h00000124;
reset = 1'b0;
P_Trace_Instruction = 32'hFA61000C;
P_Trace_Valid_Instr = 1'b1;
clk = 1'b1;
sel = 1'b0;
in_addr = 4'b0000;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000180;
reset = 1'b0;
P_Trace_Instruction = 32'h20E00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000184;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F41508;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000188;
reset = 1'b0;
P_Trace_Instruction = 32'h20A00000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000188;
reset = 1'b0;
P_Trace_Instruction = 32'h20A00000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000168C;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFE4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001690;
reset = 1'b0;
P_Trace_Instruction = 32'hFA610018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001694;
reset = 1'b0;
P_Trace_Instruction = 32'h12610000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001698;
reset = 1'b0;
P_Trace_Instruction = 32'hF8130004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000169C;
reset = 1'b0;
P_Trace_Instruction = 32'h30603590;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016A0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016A4;
reset = 1'b0;
P_Trace_Instruction = 32'h306046D0;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016A8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8130004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B0;
reset = 1'b0;
P_Trace_Instruction = 32'hB8000284;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C4;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016C8;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016CC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016D8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E0;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016E8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016EC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F4;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016F8;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000016FC;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001700;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001704;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001708;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000170C;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001710;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001714;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001718;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000171C;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001720;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001724;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001728;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000172C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001730;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001734;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001738;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000173C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001740;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001744;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001748;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000174C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001750;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001754;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001758;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000175C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001760;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001764;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001768;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000176C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001770;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001774;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001778;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000177C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001780;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001784;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001788;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000178C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001790;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001794;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001798;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000179C;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A0;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A4;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017A8;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017AC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B0;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B4;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017B8;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017BC;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C0;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017C8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017CC;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017D8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017DC;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E0;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017E8;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017EC;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F4;
reset = 1'b0;
P_Trace_Instruction = 32'h30630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000017FC;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001800;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001804;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001808;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000180C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001810;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001814;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001818;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000181C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001820;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001824;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001828;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000182C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001830;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001834;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001838;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000183C;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001840;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001844;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001848;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000184C;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001850;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001854;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001858;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000185C;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001860;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001864;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001868;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000186C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001870;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001874;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001878;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000187C;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001880;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001884;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001888;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000188C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001890;
reset = 1'b0;
P_Trace_Instruction = 32'h3063000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001894;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001898;
reset = 1'b0;
P_Trace_Instruction = 32'h88641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000189C;
reset = 1'b0;
P_Trace_Instruction = 32'hF873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A4;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018A8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018AC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018B8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018BC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018C8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018CC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018D8;
reset = 1'b0;
P_Trace_Instruction = 32'hA46300FF;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018DC;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E0;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E4;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018E8;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018EC;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F0;
reset = 1'b0;
P_Trace_Instruction = 32'hE873000C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F4;
reset = 1'b0;
P_Trace_Instruction = 32'h64630018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018F8;
reset = 1'b0;
P_Trace_Instruction = 32'hE0633490;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000018FC;
reset = 1'b0;
P_Trace_Instruction = 32'h10830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001900;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001904;
reset = 1'b0;
P_Trace_Instruction = 32'h10632000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001908;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000190C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8930004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001910;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001914;
reset = 1'b0;
P_Trace_Instruction = 32'h10641800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001918;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000191C;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001920;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001924;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001928;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730010;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000192C;
reset = 1'b0;
P_Trace_Instruction = 32'h30630010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001930;
reset = 1'b0;
P_Trace_Instruction = 32'hF8730010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001934;
reset = 1'b0;
P_Trace_Instruction = 32'hE8730014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001938;
reset = 1'b0;
P_Trace_Instruction = 32'hE8630000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000193C;
reset = 1'b0;
P_Trace_Instruction = 32'hBC23FD78;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001940;
reset = 1'b0;
P_Trace_Instruction = 32'h10600000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001944;
reset = 1'b0;
P_Trace_Instruction = 32'h10330000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001948;
reset = 1'b0;
P_Trace_Instruction = 32'hEA610018;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000194C;
reset = 1'b0;
P_Trace_Instruction = 32'h3021001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001950;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00001954;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00001954;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000018C;
reset = 1'b0;
P_Trace_Instruction = 32'h32630000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000190;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F432B4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000194;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000194;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00003444;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFF8;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00003448;
reset = 1'b0;
P_Trace_Instruction = 32'hD9E00800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000344C;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F4CC24;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00003450;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00003450;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000070;
reset = 1'b0;
P_Trace_Instruction = 32'hE06046B0;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000074;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFE4;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000074;
reset = 1'b0;
P_Trace_Instruction = 32'h3021FFE4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000078;
reset = 1'b0;
P_Trace_Instruction = 32'hBE03001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h0000007C;
reset = 1'b0;
P_Trace_Instruction = 32'hF9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000007C;
reset = 1'b0;
P_Trace_Instruction = 32'hF9E10000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000094;
reset = 1'b0;
P_Trace_Instruction = 32'hE8603488;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000094;
reset = 1'b0;
P_Trace_Instruction = 32'hE8603488;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000094;
reset = 1'b0;
P_Trace_Instruction = 32'hE8603488;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000098;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000098;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000098;
reset = 1'b0;
P_Trace_Instruction = 32'hE8830000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000009C;
reset = 1'b0;
P_Trace_Instruction = 32'hBE24FFEC;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000A0;
reset = 1'b0;
P_Trace_Instruction = 32'h30630004;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000A4;
reset = 1'b0;
P_Trace_Instruction = 32'hB0000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000A8;
reset = 1'b0;
P_Trace_Instruction = 32'h30600000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000AC;
reset = 1'b0;
P_Trace_Instruction = 32'hBC030010;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000000B0;
reset = 1'b0;
P_Trace_Instruction = 32'h30A046A4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000B0;
reset = 1'b0;
P_Trace_Instruction = 32'h30A046A4;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000BC;
reset = 1'b0;
P_Trace_Instruction = 32'h30600001;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C0;
reset = 1'b0;
P_Trace_Instruction = 32'hF06046B0;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE9E10000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C4;
reset = 1'b0;
P_Trace_Instruction = 32'hE9E10000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000C8;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000000CC;
reset = 1'b0;
P_Trace_Instruction = 32'h3021001C;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000000CC;
reset = 1'b0;
P_Trace_Instruction = 32'h3021001C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00003454;
reset = 1'b0;
P_Trace_Instruction = 32'hC9E00800;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00003454;
reset = 1'b0;
P_Trace_Instruction = 32'hC9E00800;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00003454;
reset = 1'b0;
P_Trace_Instruction = 32'hC9E00800;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00003458;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h0000345C;
reset = 1'b0;
P_Trace_Instruction = 32'h30210008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000345C;
reset = 1'b0;
P_Trace_Instruction = 32'h30210008;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000198;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F42F34;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h0000019C;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h0000019C;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000030CC;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000030D0;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000030D0;
reset = 1'b0;
P_Trace_Instruction = 32'h80000000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001A0;
reset = 1'b0;
P_Trace_Instruction = 32'hC9E10000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001A4;
reset = 1'b0;
P_Trace_Instruction = 32'h30730000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001A4;
reset = 1'b0;
P_Trace_Instruction = 32'h30730000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001A8;
reset = 1'b0;
P_Trace_Instruction = 32'hB60F0008;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h000001AC;
reset = 1'b0;
P_Trace_Instruction = 32'h20210014;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000001AC;
reset = 1'b0;
P_Trace_Instruction = 32'h20210014;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000064;
reset = 1'b0;
P_Trace_Instruction = 32'hB9F43160;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b1;
#20 P_Trace_PC = 32'h00000068;
reset = 1'b0;
P_Trace_Instruction = 32'h30A30000;
P_Trace_Valid_Instr = 1'b1;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h00000068;
reset = 1'b0;
P_Trace_Instruction = 32'h30A30000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000031C4;
reset = 1'b0;
P_Trace_Instruction = 32'hBA0C0018;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000031C4;
reset = 1'b0;
P_Trace_Instruction = 32'h10C00000;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000031C4;
reset = 1'b0;
P_Trace_Instruction = 32'hFA61001C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000031C4;
reset = 1'b0;
P_Trace_Instruction = 32'hFA61001C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000031C4;
reset = 1'b0;
P_Trace_Instruction = 32'hFA61001C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000031C4;
reset = 1'b0;
P_Trace_Instruction = 32'hFA61001C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;
#20 P_Trace_PC = 32'h000031C4;
reset = 1'b0;
P_Trace_Instruction = 32'hFA61001C;
P_Trace_Valid_Instr = 1'b0;
P_Trace_Jump_Taken = 1'b0;








//$display("ram_out=%h",uut.ram_out);
    $finish;
end

always
#10 clk=~clk;



	
      
endmodule