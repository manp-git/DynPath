`timescale 1ns / 1ps


module PDIL_PSPIC(
input clk,
input reset,
//input st4,
input st7,
input st8,
input l,
input f,
//input call,
//input loop_exit,// substuted with its expression by below two
input loop_det,
input P_Trace_Jump_Taken,
input ret,
input [4:0] match_addr,
//input code_end,
//input [4:0] f2, // delayed from f1
//input reg [4:0] f,
output reg [4:0] f2,f1,//depth of path =20, so 5 bit 
output [5:0] data_out,
output reg [19:0] flag_reg,//depth of path =20

output [4:0] next_free_location,//depth of path =20, so 5 bit 
//output reg path_return_mode, path_entry_mode,
//output reg [5:0] temp_size

output [31:0] pcam_out0,
output [31:0] pcam_out1,
output [31:0] pcam_out2,
output [31:0] pcam_out3,
output [31:0] pcam_out4,
output [31:0] pcam_out5,
output [31:0] pcam_out6,
output [31:0] pcam_out7,
output [31:0] pcam_out8,
output [31:0] pcam_out9,
output [31:0] pcam_out10,
output [31:0] pcam_out11,
output [31:0] pcam_out12,
output [31:0] pcam_out13,
output [31:0] pcam_out14,
output [31:0] pcam_out15,
output [31:0] pcam_out16,
output [31:0] pcam_out17,
output [31:0] pcam_out18,
output [31:0] pcam_out19,
output [31:0] pcam_out20,
output [31:0] pcam_out21,
output [31:0] pcam_out22,
output [31:0] pcam_out23,
output [31:0] pcam_out24,
output [31:0] pcam_out25,
output [31:0] pcam_out26,
output [31:0] pcam_out27,
output [31:0] pcam_out28,
output [31:0] pcam_out29,
output [31:0] pcam_out30,
output [31:0] pcam_out31,

output [7:0] hit_out0,
output [7:0] hit_out1,
output [7:0] hit_out2,
output [7:0] hit_out3,
output [7:0] hit_out4,
output [7:0] hit_out5,
output [7:0] hit_out6,
output [7:0] hit_out7,
output [7:0] hit_out8,
output [7:0] hit_out9,
output [7:0] hit_out10,
output [7:0] hit_out11,
output [7:0] hit_out12,
output [7:0] hit_out13,
output [7:0] hit_out14,
output [7:0] hit_out15,
output [7:0] hit_out16,
output [7:0] hit_out17,
output [7:0] hit_out18,
output [7:0] hit_out19,
output [7:0] hit_out20,
output [7:0] hit_out21,
output [7:0] hit_out22,
output [7:0] hit_out23,
output [7:0] hit_out24,
output [7:0] hit_out25,
output [7:0] hit_out26,
output [7:0] hit_out27,
output [7:0] hit_out28,
output [7:0] hit_out29,
output [7:0] hit_out30,
output [7:0] hit_out31,

output [255:0] PSPIC0,
output [255:0] PSPIC1,
output [255:0] PSPIC2,
output [255:0] PSPIC3,
output [255:0] PSPIC4,
output [255:0] PSPIC5,
output [255:0] PSPIC6,
output [255:0] PSPIC7,
output [255:0] PSPIC8,
output [255:0] PSPIC9,
output [255:0] PSPIC10,
output [255:0] PSPIC11,
output [255:0] PSPIC12,
output [255:0] PSPIC13,
output [255:0] PSPIC14,
output [255:0] PSPIC15,
output [255:0] PSPIC16,
output [255:0] PSPIC17,
output [255:0] PSPIC18,
output [255:0] PSPIC19,
output [255:0] PSPIC20,
output [255:0] PSPIC21,
output [255:0] PSPIC22,
output [255:0] PSPIC23,
output [255:0] PSPIC24,
output [255:0] PSPIC25,
output [255:0] PSPIC26,
output [255:0] PSPIC27,
output [255:0] PSPIC28,
output [255:0] PSPIC29,
output [255:0] PSPIC30,
output [255:0] PSPIC31
//output [255:0] PSPIC32

    );
	 
wire temp_switch_pulse;	 
wire temp_length;
 /*(* keep = "true" *)*/ reg [4:0] flag_addr [23:0]; //max. depth of path=20 //cam tag=6bits
 /*(* keep = "true" *) */reg [4:0] path_temp [23:0]; //max. depth of path=20
 /*(* keep = "true" *)*/ reg [4:0] path_temp_d1 [23:0]; //max. depth of path=20


 /*(* keep = "true" *) */reg [7:0] ps_invc [31:0]; //max. no. of process profiler supports
 /*(* keep = "true" *)*/ reg [7:0] ps_invc_temp [31:0]; //max. no. of process profiler supports

 //(* keep = "true" *)
  //reg [255:0] PSPIC [31:0];
 (* ram_style = "distributed" *) reg [255:0] PSPIC [31:0];
reg [4:0] temp_size;//temp size for CAM folding condition
reg [4:0] next_free_loc;//depth of path =20, so 5 bit 
reg [4:0] branching_pointer_old, branching_pointer_new;//depth of path =20, so 5 bit 

reg temp_switch, temp_switch_d1;
reg st7_d1;
reg st7_d2;

integer i,j,k,m,n,h,w;//loop index
wire [1:0] length_path;

always@(posedge clk)
begin
    if(reset)
    begin
        st7_d1 <= 1'b0;

        end
    else
    begin
  // st6_d1<=st6;
        st7_d1 <=  st7;

end
end
always@(posedge clk)
begin
    if(reset)
    begin
  //  st6_d2<=1'b0;
        st7_d2 <= 1'b0;

        end
    else
    begin
   // st6_d2<=st6_d1;
        st7_d2 <=  st7_d1;

end
end





/* --------------------------------------- TRACKING PURPOSE --------------------------------------*/
always @ (posedge clk)
begin
if(reset) begin

  next_free_loc <= 5'b0;
  //temp_to_cam<=1'b0;
//  path_temp_sel<= 1'b0;
  temp_switch = 1'b1;
  temp_size<=5'b0;
  f2<=5'b00000; 
  f1<=5'b00000;
  flag_reg<=40'b0;
  branching_pointer_old<=5'b0; //to consider for current path
  branching_pointer_new<=5'b0; // to consider for next path
  i=0;
  j=0;
  k=0;
  m=0;
  n=0;
  h=0;
  w=0;
  
  flag_addr[0] <= 5'b0;
  flag_addr[1] <= 5'b0;
  flag_addr[2] <= 5'b0;
  flag_addr[3] <= 5'b0;
  flag_addr[4] <= 5'b0;
  flag_addr[5] <= 5'b0;
  flag_addr[6] <= 5'b0;
  flag_addr[7] <= 5'b0;
  flag_addr[8] <= 5'b0;
  flag_addr[9] <= 5'b0;
  flag_addr[10] <=5'b0;
  flag_addr[11] <= 5'b0;
  flag_addr[12] <= 5'b0;
  flag_addr[13] <= 5'b0;
  flag_addr[14] <= 5'b0;
  flag_addr[15] <= 5'b0;
  flag_addr[16] <= 5'b0;
  flag_addr[17] <= 5'b0;
  flag_addr[18] <= 5'b0;
  flag_addr[19] <= 5'b0;
  flag_addr[20] <= 5'b0;
  flag_addr[21] <= 5'b0;
  flag_addr[22] <= 5'b0;
  flag_addr[23] <= 5'b0;
  
   path_temp[0] <= 5'b0;
   path_temp[1] <= 5'b0;
   path_temp[2] <= 5'b0;
   path_temp[3] <= 5'b0;
   path_temp[4] <= 5'b0;
   path_temp[5] <= 5'b0;
   path_temp[6] <= 5'b0;
   path_temp[7] <= 5'b0;
   path_temp[8] <= 5'b0;
   path_temp[9] <= 5'b0;
   path_temp[10] <= 5'b0;
   path_temp[11] <= 5'b0;
   path_temp[12] <= 5'b0;
   path_temp[13] <= 5'b0;
   path_temp[14] <= 5'b0;
   path_temp[15] <= 5'b0;
   path_temp[16] <= 5'b0;
   path_temp[17] <= 5'b0;
   path_temp[18] <= 5'b0;
   path_temp[19] <= 5'b0; 
   path_temp[20] <= 5'b0;
   path_temp[21] <= 5'b0;
   path_temp[22] <= 5'b0;
   path_temp[23] <= 5'b0;
   
  ps_invc[0] <= 8'b0;
  ps_invc[1] <= 8'b0;
  ps_invc[2] <= 8'b0;
  ps_invc[3] <= 8'b0;
  ps_invc[4] <= 8'b0;
  ps_invc[5] <= 8'b0;
  ps_invc[6] <= 8'b0;
  ps_invc[7] <= 8'b0;
  ps_invc[8] <= 8'b0;
  ps_invc[9] <= 8'b0;
  ps_invc[10] <=8'b0;
  ps_invc[11] <= 8'b0;
  ps_invc[12] <= 8'b0;
  ps_invc[13] <= 8'b0;
  ps_invc[14] <= 8'b0;
  ps_invc[15] <= 8'b0;
  ps_invc[16] <= 8'b0;
  ps_invc[17] <= 8'b0;
  ps_invc[18] <= 8'b0;
  ps_invc[19] <= 8'b0;
  ps_invc[20] <= 8'b0;
  ps_invc[21] <= 8'b0;
  ps_invc[22] <= 8'b0;
  ps_invc[23] <= 8'b0;
 /* ps_invc[24] <= 8'b0;
  ps_invc[25] <= 8'b0;
  ps_invc[26] <= 8'b0;
  ps_invc[27] <= 8'b0;
  ps_invc[28] <= 8'b0;
  ps_invc[29] <= 8'b0;
  ps_invc[30] <=8'b0;
  ps_invc[31] <= 8'b0;*/
 
 
  ps_invc_temp[0] <= 8'b0;
  ps_invc_temp[1] <= 8'b0;
  ps_invc_temp[2] <= 8'b0;
  ps_invc_temp[3] <= 8'b0;
  ps_invc_temp[4] <= 8'b0;
  ps_invc_temp[5] <= 8'b0;
  ps_invc_temp[6] <= 8'b0;
  ps_invc_temp[7] <= 8'b0;
  ps_invc_temp[8] <= 8'b0;
  ps_invc_temp[9] <= 8'b0;
  ps_invc_temp[10] <=8'b0;
  ps_invc_temp[11] <= 8'b0;
  ps_invc_temp[12] <= 8'b0;
  ps_invc_temp[13] <= 8'b0;
  ps_invc_temp[14] <= 8'b0;
  ps_invc_temp[15] <= 8'b0;
  ps_invc_temp[16] <= 8'b0;
  ps_invc_temp[17] <= 8'b0;
  ps_invc_temp[18] <= 8'b0;
  ps_invc_temp[19] <= 8'b0;
  ps_invc_temp[20] <= 8'b0;
  ps_invc_temp[21] <= 8'b0;
  ps_invc_temp[22] <= 8'b0;
  ps_invc_temp[23] <= 8'b0;
/*  ps_invc_temp[24] <= 8'b0;
  ps_invc_temp[25] <= 8'b0;
  ps_invc_temp[26] <= 8'b0;
  ps_invc_temp[27] <= 8'b0;
  ps_invc_temp[28] <= 8'b0;
  ps_invc_temp[29] <= 8'b0;
  ps_invc_temp[30] <=8'b0;
  ps_invc_temp[31] <= 8'b0;*/
 
   

   end
 
	
	//ENTRY 
else if((st7 &l)|| (st7_d2 &f))  // from st7_d1 &l in questa
 begin
   
 //CASE-1  
	 if((f2==5'b00000) && (f1==5'b00000)) 
         begin 
	       //  f1<=next_free_loc;//f2
	         f1<=f2;//7-1-2021
	       //  flag_addr[next_free_loc]<= match_addr; //f2
	         flag_addr[f2]<= match_addr; //7-1-2021
	      //   f2<=next_free_loc+1;//f2+6'b000001; 
	         ps_invc[f2] <= ps_invc[f2]+1'b1;
	         f2<=f2+5'b00001;//7-1-2021; 
	     //    flag_reg[next_free_loc]<=1'b1; //17-12-2020 for hit2 //flag_reg[f1]<=1'b1;...........TEST HIT 1 AGAIN AND ANALYSE
	         flag_reg[f1]<=1'b1;//7-1-2021;
	         //  path_return_mode<=1'b0;      // reset path pointer has started
             //	path_entry_mode <= 1'b1;
		   //  next_free_loc<= next_free_loc+1; //26-11-2020  
		     next_free_loc<= 1'b1; //7-1-2021
	     end
	     
//CASE-2    //Detect change required in Current position and for the forward direction
	  else if (flag_addr[f2-1]!=match_addr) 
	      begin 
	         if (f2==next_free_loc) //-> no matchrequired, just fill AS USUAL
	             begin
	                f1<=f2;
	                flag_addr[next_free_loc]<=match_addr;
	                ps_invc[next_free_loc] <= ps_invc[next_free_loc]+1'b1;
	                
 	                f2<=f2+5'b00001;
	                flag_reg[f1+1]<=1'b1;
	                next_free_loc<= next_free_loc+1;
	             end
	    

	         else if (f2<next_free_loc) // -> match required
	             begin
	                if (flag_addr[f2]==match_addr) //equal then continue- path retracing itself or loop
	                    begin
	                       f1<=f2;//26-11-2020
	                      f2<=f2+5'b00001;
	                       ps_invc[f2] <= ps_invc[f2]+1'b1;
	                       flag_reg[f1+1]<=1'b1;//26-11-2020
	                       next_free_loc<= next_free_loc;
	                    end
	  //culprit - 1st ques why f2<next_loc             
	                else if (flag_addr[f2]!=match_addr)//) || (f2==6'b0 && (ret )))// -> different means tempswitch //branchchange
	                //copy parent path
	                    begin
	                        branching_pointer_old<=branching_pointer_new;
	                        branching_pointer_new <= f2;
	                        for(k=0; k<24; k=k+1) begin
	                          if(k<20) begin // parent path copy
	                          path_temp[k]<=flag_addr[k]; //end
	                          ps_invc_temp[k]<= ps_invc[k]; end
	                          if(k==f2) begin // replace with new addr
	                          flag_addr[k]<= match_addr;// end
	                          ps_invc[k]<=1; end
	                          if(k>f2) begin // to replace all existing values with all zeroes
	                          flag_addr[k]<=0; //end
	                         ps_invc[k]<=0; end
	                        end                 
	                                       
	                    /*copy data to temp path
	                    put a generate loop - for index>f2=0
	                    f2=nw
	                    rest as it is*/
	                       f1<=f2;//26-11-2020
	                       f2<=f2+5'b00001;
	                       flag_reg[f1+1]<=1'b1;//26-11-2020
	                       temp_switch<=~temp_switch;//yet to decide
	                       temp_size<=next_free_loc;//yet to decide
	                       next_free_loc<=f2+1;
	                       
	                   //    length_path<=(3<=next_free_loc<=5)?2'b01:(1<=next_free_loc<=2)?2'b10:2'b00;
	                       
	                    //   f1<=0;
	                  //     f2<=0;
	                    end 
	              end
	          else;
           end	       
  end


	 
else if (st8 & (ret | (loop_det & !P_Trace_Jump_Taken)))//both logical and arith and-or are fine
//(st8 && (ret || loop_exit)) with loop_exit- simulator was getting loop_exit-1 not at correct instance, though it was 1 in that clock cycle..
//i.e. loop_det was 1 but loop exit was 0 at initial instance// it was all issue wrt simulator sequencing, with description inside flag_arrd of loop exit - it works fine
	   begin 
	      if(f2==5'b00001) begin // chks old value of f //Takes care of last ret/exit form user code
	      //done to take care of 1-2 = 1f issue in f1 variable
	         f1<= f2-5'b00001; 
	// COPY ENTIRE PATH WHEN EXIT TO MAIN        

	         for(n=0; n<24; n=n+1) 
	           begin
	             path_temp[n]<=flag_addr[n]; 
	           end

	         temp_switch<=~temp_switch;//yet to decide
	         temp_size<=next_free_loc;//yet to decide
	         next_free_loc<=0;
	         
	       //  length_path<=(3<=next_free_loc<=5)?2'b01:(1<=next_free_loc<=2)?2'b10:2'b00;
	      end
	         
	      else begin
	           f1<= f2-5'b00010; 
	         	     // next_free_loc<= next_free_loc;
	           end  
	   
	      f2<=f2-5'b00001; 
	      flag_reg[f1]<=1'b0;
	         
	   end //end st8
	          //nonblocking assignments evaluated first updated later
	         // if blocking behaves full sequentially, then f1<= f-5'b00001;
	         
else;

end

/* --------------------------------------- MATCHING PURPOSE --------------------------------------*/
//path switch indication to matching forward
always@(posedge clk)
begin
    if(reset)
        temp_switch_d1 <= 1'b0;
    else temp_switch_d1 <= temp_switch;
end

assign temp_switch_pulse = (temp_switch ^ temp_switch_d1);

wire [119:0] path_temp_combined;
//coverts vertical pathtemp reg to one horizontal vector for matching purpose
assign path_temp_combined = {path_temp[19],path_temp[18],path_temp[17],path_temp[16],path_temp[15],path_temp[14],path_temp[13],path_temp[12],path_temp[11],path_temp[10],path_temp[9],path_temp[8],path_temp[7],path_temp[6],path_temp[5],path_temp[4],path_temp[3],path_temp[2],path_temp[1],path_temp[0]};

// SEPARATION INTO dual path temp reg for matching purpose
reg [119:0] path_temp0,path_temp1;
//reg [99:0] path_temp0,path_temp1;
always@(*)
begin
path_temp0<=(reset)?120'b0:(temp_switch_pulse & temp_switch)?path_temp_combined:path_temp0;
path_temp1<=(reset)?120'b0:(temp_switch_pulse & (!temp_switch))?path_temp_combined:path_temp1;
end

/***********common_TPR / counter for verification purpose only****************/
reg [119:0] common_TPR;
//reg [89:0] common_TPR;
//reg [29:0] test_count0, test_count1, test_count2, test_count3, test_count4, test_count5, test_count6, test_count7, test_count8, test_count9, test_count10;

always@(posedge clk)
begin
if (reset)
begin
common_TPR<= 120'b0;

end

else if(temp_switch_pulse)
begin
// hardware pupose - common_TPR<= temp_switch ? path_temp0:path_temp1;//(temp_switch & path_temp0);// | ((~temp_switch) && path_temp1);

/***********counter for verification purpose only****************/
common_TPR= temp_switch ? path_temp0:path_temp1;//(temp_switch & path_temp0);// | ((~temp_switch) && path_temp1);

/****************************/
end
end
/****************************/

assign data_out = flag_addr[f1];
assign next_free_location = next_free_loc;

//assign length_path=((temp_size>=16)&&(temp_size<=20))?2'b11:((temp_size>=11)&&(temp_size<=15))?2'b10:((temp_size>=6)&&(temp_size<=10))?2'b01:2'b00;
assign length_path=((temp_size>=19)&&(temp_size<=24))?2'b11:((temp_size>=13)&&(temp_size<=18))?2'b10:((temp_size>=7)&&(temp_size<=12))?2'b01:2'b00;
/////////////////////////////////////

reg [3:0] cam_state, next_state;
reg [4:0] read_addr, path_addr,path_count,p;
reg [119:0] MatchReg;
reg [31:0] cam [31:0];
reg A,B,C,D;
reg [5:0] wr_addr; // 1 extra bit so as to not overlap with 0 on a safer side
reg hit_wren;


parameter S0 = 4'b0000;
parameter S1 = 4'b0001;
parameter S2 = 4'b0010;
parameter S3 = 4'b0011;
parameter S4 = 4'b0100;
parameter S5 = 4'b0101;
parameter S6 = 4'b0110;
parameter S7 = 4'b0111;

 
always @(posedge clk)
begin
	if(reset)    // not rst_int 
	cam_state <= S0;
	else
	cam_state <= next_state;
end

always@(posedge clk)
begin
for (m=0;m<24;m=m+1)
begin
if (reset)
begin
path_temp_d1[m]<=0;
//path_temp_d2[m]<=0;
end
else begin
path_temp_d1[m]<=path_temp[m];
//path_temp_d2[m]<=path_temp_d1[m];
end
end
end

 //cam0 filling pending
 always@(*)
 //always@(posedge clk) - synth error
 begin
    //next_state=S_INIT;
    case(cam_state)
    
        S0://reset and state
            begin
                read_addr=0;
                path_addr=0;
                MatchReg=0;
                wr_addr=0;
                A=0;
                B=0;
                C=0;
                D=0;
                cam[0]=0;
                cam[1]=0;
                cam[2]=0;
                cam[3]=0;
                cam[4]=0;
                cam[5]=0;    
                cam[6]=0;
                cam[7]=0;
                cam[8]=0;
                cam[9]=0;
                cam[10]=0;
                cam[11]=0;
                cam[12]=0;
                cam[13]=0;
                cam[14]=0;
                cam[15]=0;    
                cam[16]=0;
                cam[17]=0;
                cam[18]=0;
                cam[19]=0;
                cam[20]=0;
                cam[21]=0;
                cam[22]=0;
                cam[23]=0;
                cam[24]=0;
                cam[25]=0;    
                cam[26]=0;
                cam[27]=0;
                cam[28]=0;
                cam[29]=0;
                cam[30]=0;
                cam[31]=0;
                path_count=0;
                p=0;                           
                next_state=S1;
                hit_wren = 1'b0;

            end
                
        S1: //WAIT
            begin
                hit_wren = 1'b0;
                read_addr=0;
                p=1;// as used only in case of cam not empty which also means atleast 1 path already in it, so p starts from 1 and path_count also is atleast 1 and S2 executes atleast once post this  which means all are fine parallely
                if (temp_switch_pulse & cam[0][0]==0)//empty cam
                next_state= S4;//empty cam fill state
                else if (temp_switch_pulse & (!cam[0][0]==0))
                next_state= S2; //load match reg state
            end
        S2: //read addr is required to be 0 after S0, updated as per closing after 
            begin //LOAD MATCH REG
                A= cam[read_addr][0];
                B= cam[read_addr+1][0];
                C= cam[read_addr+2][0];
                D= cam[read_addr+3][0];
                MatchReg[29:0]=(A)?cam[read_addr][31:2]:30'b0;  //ACTUALLY DONT NEED TO WRITE AS A HERE, ANYHOW FOR A=1 IS WHEN FILL MATCH REG UNLIKE BELOW WHR FILL ON 0;
                MatchReg[59:30]=(B)?30'b0:cam[read_addr+1][31:2];
                MatchReg[89:60]=(B|C)?30'b0:cam[read_addr+2][31:2]; // corrected from + to | as + will add not required result overflows and result of B+C is 10 and not 1
                MatchReg[119:90]=(B|C|D)?30'b0:cam[read_addr+3][31:2];
                                                  
                next_state=S3;
                hit_wren = 1'b0;
             end
                         
         S3://match state
             begin

                if (MatchReg==common_TPR)
                //next_state= S4;
                begin  path_addr=read_addr;
                hit_wren = 1'b1;
                next_state=S1; 
	               
   		 
          
                end
 
                
                else
                    begin
                        next_state= (p<path_count)?S2:S5; //when not match proceed further
                     //   READ_ADDR MANIP USING EXISTING A,B,C,D VALUES
                    // SO AS TO FIND NEXT A=1 POSITION.
                        read_addr= (p<path_count)?(A&B)?read_addr+1:(A&(~B)&C)?read_addr+2:(A&(~B)&(~C)&D)?read_addr+3:(A&(~B)&(~C)&(~D))?read_addr+4:0:read_addr; // could be read_addr:read_addr also?
                        p=p+1;//whr put doesnt matter 
                        
                    //    LOOPING HERE BETWEEN s1&s2 - WHAT IF NO MATCH-- Added S4 ANDPASS ON READ ADDR FOR TO GET STORED IN S4
                        
                    end
                end
         S4:// cam write when cam empty
            begin
                path_addr=5'b0;
                hit_wren = 1'b1;
                //read_addr=5'b0;////////no zero put logic here
            //    wr_en=1; //////no need to do write en high- just put write logic directly as fsm is coordinating already, no separate block required
                next_state=S1;    

                cam[wr_addr]= {common_TPR[29:0],2'b01};
                cam[wr_addr+1]= (length_path>=2)? {common_TPR[59:30],2'b00}:32'b0;
                cam[wr_addr+2]= (length_path>=3)? {common_TPR[89:60],2'b00}:32'b0;
                cam[wr_addr+3]= (length_path>=4)? {common_TPR[119:90],2'b00}:32'b0;
                path_count=path_count+1;
                
      

                wr_addr= wr_addr+length_path+1;// as path length is 0 to 3
         //       wr_addr=last filled based on length path;        -- follow read_addr logic                      
                             
            end
            
         S5: //cam write when not empty
            begin
                path_addr= read_addr+l; // 20-mar-2021 corrected from read_addr .. WHY+1, should be based on length of previous path 28-Mar-2021
              //  wr_en=1;
                next_state=S1;
                hit_wren = 1'b1;
             
                cam[wr_addr]= {common_TPR[29:0],2'b01};
                cam[wr_addr+1]= (length_path>=2)? {common_TPR[59:30],2'b00}:32'b0;
                cam[wr_addr+2]= (length_path>=3)? {common_TPR[89:60],2'b00}:32'b0;
                cam[wr_addr+3]= (length_path>=4)? {common_TPR[119:90],2'b00}:32'b0;
                path_count=path_count+1;
                wr_addr= wr_addr+length_path+1;// as path length is 0 to 3
        //        wr_addr=last filled based on length path;        -- follow read_addr logic 
		       
 
                     
             end
                       
          	   default: next_state = S0;
		
		endcase
          
    end


wire hit_wr_en;
reg [4:0] path_addr_d1;

always@(posedge clk)
begin
    if(reset)
    begin
        path_addr_d1<=5'b0;
        end
    else
    begin
        path_addr_d1<=path_addr;
end
end

assign hit_wr_en = hit_wren; 

always @ (posedge clk)
begin
if (reset)
begin
     for (h=0;h<32;h=h+1)
       begin
           PSPIC[h]=0;
       end 
end
else if (hit_wr_en)
begin
              case(path_addr_d1)
                5'd0 : begin
                    PSPIC[path_temp_d1[0]][7:0]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][7:0]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][7:0];
                    PSPIC[path_temp_d1[1]][7:0]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][7:0]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][7:0];
                    PSPIC[path_temp_d1[2]][7:0]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][7:0]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][7:0];
                    PSPIC[path_temp_d1[3]][7:0]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][7:0]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][7:0];
                    PSPIC[path_temp_d1[4]][7:0]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][7:0]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][7:0];
                    PSPIC[path_temp_d1[5]][7:0]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][7:0]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][7:0];
                    PSPIC[path_temp_d1[6]][7:0]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][7:0]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][7:0];
                    PSPIC[path_temp_d1[7]][7:0]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][7:0]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][7:0];
                    PSPIC[path_temp_d1[8]][7:0]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][7:0]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][7:0];
                    PSPIC[path_temp_d1[9]][7:0]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][7:0]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][7:0];
                    PSPIC[path_temp_d1[10]][7:0]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][7:0]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][7:0];
                    PSPIC[path_temp_d1[11]][7:0]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][7:0]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][7:0];
                    PSPIC[path_temp_d1[12]][7:0]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][7:0]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][7:0];
                    PSPIC[path_temp_d1[13]][7:0]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][7:0]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][7:0];
                    PSPIC[path_temp_d1[14]][7:0]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][7:0]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][7:0];
                    PSPIC[path_temp_d1[15]][7:0]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][7:0]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][7:0];
                    PSPIC[path_temp_d1[16]][7:0]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][7:0]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][7:0];
                    PSPIC[path_temp_d1[17]][7:0]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][7:0]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][7:0];
                    PSPIC[path_temp_d1[18]][7:0]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][7:0]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][7:0];
                    PSPIC[path_temp_d1[19]][7:0]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][7:0]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][7:0];
                    PSPIC[path_temp_d1[20]][7:0]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][7:0]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][7:0];
                    PSPIC[path_temp_d1[21]][7:0]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][7:0]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][7:0];
                    PSPIC[path_temp_d1[22]][7:0]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][7:0]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][7:0];
                    PSPIC[path_temp_d1[23]][7:0]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][7:0]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][7:0];             
                     end
                     
              /*   5'd0 : begin
                    PSPIC[path_temp_d1[0]][7:0]<=(0>=branching_pointer_old)?(ps_invc_temp[0]):PSPIC[path_temp_d1[0]][7:0];
                    PSPIC[path_temp_d1[1]][7:0]<=(1>=branching_pointer_old)?(ps_invc_temp[1]):PSPIC[path_temp_d1[1]][7:0];
                    PSPIC[path_temp_d1[2]][7:0]<=(2>=branching_pointer_old)?(ps_invc_temp[2]):PSPIC[path_temp_d1[2]][7:0];
                    PSPIC[path_temp_d1[3]][7:0]<=(3>=branching_pointer_old)?(ps_invc_temp[3]):PSPIC[path_temp_d1[3]][7:0];
                    PSPIC[path_temp_d1[4]][7:0]<=(4>=branching_pointer_old)?(ps_invc_temp[4]):PSPIC[path_temp_d1[4]][7:0];
                    PSPIC[path_temp_d1[5]][7:0]<=(5>=branching_pointer_old)?(ps_invc_temp[5]):PSPIC[path_temp_d1[5]][7:0];
                    PSPIC[path_temp_d1[6]][7:0]<=(6>=branching_pointer_old)?(ps_invc_temp[6]):PSPIC[path_temp_d1[6]][7:0];
                    PSPIC[path_temp_d1[7]][7:0]<=(7>=branching_pointer_old)?(ps_invc_temp[7]):PSPIC[path_temp_d1[7]][7:0];
                    PSPIC[path_temp_d1[8]][7:0]<=(8>=branching_pointer_old)?(ps_invc_temp[8]):PSPIC[path_temp_d1[8]][7:0];
                    PSPIC[path_temp_d1[9]][7:0]<=(9>=branching_pointer_old)?(ps_invc_temp[9]):PSPIC[path_temp_d1[9]][7:0];
                    PSPIC[path_temp_d1[10]][7:0]<=(10>=branching_pointer_old)?(ps_invc_temp[10]):PSPIC[path_temp_d1[10]][7:0];
                    PSPIC[path_temp_d1[11]][7:0]<=(11>=branching_pointer_old)?(ps_invc_temp[11]):PSPIC[path_temp_d1[11]][7:0];
                    PSPIC[path_temp_d1[12]][7:0]<=(12>=branching_pointer_old)?(ps_invc_temp[12]):PSPIC[path_temp_d1[12]][7:0];
                    PSPIC[path_temp_d1[13]][7:0]<=(13>=branching_pointer_old)?(ps_invc_temp[13]):PSPIC[path_temp_d1[13]][7:0];
                    PSPIC[path_temp_d1[14]][7:0]<=(14>=branching_pointer_old)?(ps_invc_temp[14]):PSPIC[path_temp_d1[14]][7:0];
                    PSPIC[path_temp_d1[15]][7:0]<=(15>=branching_pointer_old)?(ps_invc_temp[15]):PSPIC[path_temp_d1[15]][7:0];
                    PSPIC[path_temp_d1[16]][7:0]<=(16>=branching_pointer_old)?(ps_invc_temp[16]):PSPIC[path_temp_d1[16]][7:0];
                    PSPIC[path_temp_d1[17]][7:0]<=(17>=branching_pointer_old)?(ps_invc_temp[17]):PSPIC[path_temp_d1[17]][7:0];
                    PSPIC[path_temp_d1[18]][7:0]<=(18>=branching_pointer_old)?(ps_invc_temp[18]):PSPIC[path_temp_d1[18]][7:0];
                    PSPIC[path_temp_d1[19]][7:0]<=(19>=branching_pointer_old)?(ps_invc_temp[19]):PSPIC[path_temp_d1[19]][7:0];
                    PSPIC[path_temp_d1[20]][7:0]<=(20>=branching_pointer_old)?(ps_invc_temp[20]):PSPIC[path_temp_d1[20]][7:0];
                    PSPIC[path_temp_d1[21]][7:0]<=(21>=branching_pointer_old)?(ps_invc_temp[21]):PSPIC[path_temp_d1[21]][7:0];
                    PSPIC[path_temp_d1[22]][7:0]<=(22>=branching_pointer_old)?(ps_invc_temp[22]):PSPIC[path_temp_d1[22]][7:0];
                    PSPIC[path_temp_d1[23]][7:0]<=(23==branching_pointer_old)?(ps_invc_temp[23]):PSPIC[path_temp_d1[23]][7:0];             
                     end*/
                5'd1 : begin
                    PSPIC[path_temp_d1[0]][15:8]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][15:8]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][15:8];
                    PSPIC[path_temp_d1[1]][15:8]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][15:8]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][15:8];
                    PSPIC[path_temp_d1[2]][15:8]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][15:8]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][15:8];
                    PSPIC[path_temp_d1[3]][15:8]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][15:8]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][15:8];
                    PSPIC[path_temp_d1[4]][15:8]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][15:8]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][15:8];
                    PSPIC[path_temp_d1[5]][15:8]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][15:8]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][15:8];
                    PSPIC[path_temp_d1[6]][15:8]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][15:8]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][15:8];
                    PSPIC[path_temp_d1[7]][15:8]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][15:8]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][15:8];
                    PSPIC[path_temp_d1[8]][15:8]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][15:8]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][15:8];
                    PSPIC[path_temp_d1[9]][15:8]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][15:8]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][15:8];
                    PSPIC[path_temp_d1[10]][15:8]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][15:8]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][15:8];
                    PSPIC[path_temp_d1[11]][15:8]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][15:8]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][15:8];
                    PSPIC[path_temp_d1[12]][15:8]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][15:8]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][15:8];
                    PSPIC[path_temp_d1[13]][15:8]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][15:8]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][15:8];
                    PSPIC[path_temp_d1[14]][15:8]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][15:8]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][15:8];
                    PSPIC[path_temp_d1[15]][15:8]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][15:8]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][15:8];
                    PSPIC[path_temp_d1[16]][15:8]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][15:8]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][15:8];
                    PSPIC[path_temp_d1[17]][15:8]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][15:8]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][15:8];
                    PSPIC[path_temp_d1[18]][15:8]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][15:8]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][15:8];
                    PSPIC[path_temp_d1[19]][15:8]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][15:8]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][15:8];
                    PSPIC[path_temp_d1[20]][15:8]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][15:8]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][15:8];
                    PSPIC[path_temp_d1[21]][15:8]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][15:8]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][15:8];
                    PSPIC[path_temp_d1[22]][15:8]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][15:8]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][15:8];
                    PSPIC[path_temp_d1[23]][15:8]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][15:8]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][15:8];  
                     end
                5'd2 : begin
                    PSPIC[path_temp_d1[0]][23:16]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][23:16]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][23:16];
                    PSPIC[path_temp_d1[1]][23:16]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][23:16]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][23:16];
                    PSPIC[path_temp_d1[2]][23:16]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][23:16]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][23:16];
                    PSPIC[path_temp_d1[3]][23:16]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][23:16]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][23:16];
                    PSPIC[path_temp_d1[4]][23:16]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][23:16]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][23:16];
                    PSPIC[path_temp_d1[5]][23:16]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][23:16]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][23:16];
                    PSPIC[path_temp_d1[6]][23:16]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][23:16]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][23:16];
                    PSPIC[path_temp_d1[7]][23:16]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][23:16]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][23:16];
                    PSPIC[path_temp_d1[8]][23:16]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][23:16]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][23:16];
                    PSPIC[path_temp_d1[9]][23:16]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][23:16]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][23:16];
                    PSPIC[path_temp_d1[10]][23:16]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][23:16]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][23:16];
                    PSPIC[path_temp_d1[11]][23:16]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][23:16]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][23:16];
                    PSPIC[path_temp_d1[12]][23:16]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][23:16]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][23:16];
                    PSPIC[path_temp_d1[13]][23:16]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][23:16]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][23:16];
                    PSPIC[path_temp_d1[14]][23:16]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][23:16]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][23:16];
                    PSPIC[path_temp_d1[15]][23:16]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][23:16]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][23:16];
                    PSPIC[path_temp_d1[16]][23:16]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][23:16]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][23:16];
                    PSPIC[path_temp_d1[17]][23:16]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][23:16]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][23:16];
                    PSPIC[path_temp_d1[18]][23:16]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][23:16]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][23:16];
                    PSPIC[path_temp_d1[19]][23:16]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][23:16]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][23:16];
                    PSPIC[path_temp_d1[20]][23:16]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][23:16]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][23:16];
                    PSPIC[path_temp_d1[21]][23:16]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][23:16]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][23:16];
                    PSPIC[path_temp_d1[22]][23:16]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][23:16]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][23:16];
                    PSPIC[path_temp_d1[23]][23:16]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][23:16]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][23:16];
             
                     end
                5'd3 : begin
                    PSPIC[path_temp_d1[0]][31:24]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][31:24]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][31:24];
                    PSPIC[path_temp_d1[1]][31:24]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][31:24]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][31:24];
                    PSPIC[path_temp_d1[2]][31:24]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][31:24]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][31:24];
                    PSPIC[path_temp_d1[3]][31:24]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][31:24]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][31:24];
                    PSPIC[path_temp_d1[4]][31:24]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][31:24]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][31:24];
                    PSPIC[path_temp_d1[5]][31:24]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][31:24]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][31:24];
                    PSPIC[path_temp_d1[6]][31:24]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][31:24]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][31:24];
                    PSPIC[path_temp_d1[7]][31:24]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][31:24]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][31:24];
                    PSPIC[path_temp_d1[8]][31:24]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][31:24]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][31:24];
                    PSPIC[path_temp_d1[9]][31:24]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][31:24]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][31:24];
                    PSPIC[path_temp_d1[10]][31:24]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][31:24]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][31:24];
                    PSPIC[path_temp_d1[11]][31:24]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][31:24]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][31:24];
                    PSPIC[path_temp_d1[12]][31:24]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][31:24]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][31:24];
                    PSPIC[path_temp_d1[13]][31:24]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][31:24]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][31:24];
                    PSPIC[path_temp_d1[14]][31:24]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][31:24]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][31:24];
                    PSPIC[path_temp_d1[15]][31:24]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][31:24]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][31:24];
                    PSPIC[path_temp_d1[16]][31:24]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][31:24]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][31:24];
                    PSPIC[path_temp_d1[17]][31:24]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][31:24]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][31:24];
                    PSPIC[path_temp_d1[18]][31:24]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][31:24]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][31:24];
                    PSPIC[path_temp_d1[19]][31:24]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][31:24]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][31:24];
                    PSPIC[path_temp_d1[20]][31:24]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][31:24]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][31:24];
                    PSPIC[path_temp_d1[21]][31:24]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][31:24]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][31:24];
                    PSPIC[path_temp_d1[22]][31:24]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][31:24]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][31:24];
                    PSPIC[path_temp_d1[23]][31:24]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][31:24]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][31:24];
                     end
                5'd4 : begin
                    PSPIC[path_temp_d1[0]][39:32]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][39:32]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][39:32];
                    PSPIC[path_temp_d1[1]][39:32]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][39:32]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][39:32];
                    PSPIC[path_temp_d1[2]][39:32]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][39:32]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][39:32];
                    PSPIC[path_temp_d1[3]][39:32]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][39:32]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][39:32];
                    PSPIC[path_temp_d1[4]][39:32]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][39:32]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][39:32];
                    PSPIC[path_temp_d1[5]][39:32]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][39:32]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][39:32];
                    PSPIC[path_temp_d1[6]][39:32]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][39:32]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][39:32];
                    PSPIC[path_temp_d1[7]][39:32]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][39:32]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][39:32];
                    PSPIC[path_temp_d1[8]][39:32]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][39:32]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][39:32];
                    PSPIC[path_temp_d1[9]][39:32]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][39:32]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][39:32];
                    PSPIC[path_temp_d1[10]][39:32]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][39:32]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][39:32];
                    PSPIC[path_temp_d1[11]][39:32]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][39:32]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][39:32];
                    PSPIC[path_temp_d1[12]][39:32]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][39:32]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][39:32];
                    PSPIC[path_temp_d1[13]][39:32]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][39:32]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][39:32];
                    PSPIC[path_temp_d1[14]][39:32]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][39:32]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][39:32];
                    PSPIC[path_temp_d1[15]][39:32]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][39:32]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][39:32];
                    PSPIC[path_temp_d1[16]][39:32]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][39:32]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][39:32];
                    PSPIC[path_temp_d1[17]][39:32]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][39:32]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][39:32];
                    PSPIC[path_temp_d1[18]][39:32]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][39:32]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][39:32];
                    PSPIC[path_temp_d1[19]][39:32]<=(19==branching_pointer_old)?(PSPIC[path_temp_d1[19]][39:32]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][39:32];
                    PSPIC[path_temp_d1[20]][39:32]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][39:32]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][39:32];
                    PSPIC[path_temp_d1[21]][39:32]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][39:32]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][39:32];
                    PSPIC[path_temp_d1[22]][39:32]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][39:32]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][39:32];
                    PSPIC[path_temp_d1[23]][39:32]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][39:32]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][39:32]; end
                5'd5 : begin
                    PSPIC[path_temp_d1[0]][47:40]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][47:40]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][47:40];
                    PSPIC[path_temp_d1[1]][47:40]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][47:40]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][47:40];
                    PSPIC[path_temp_d1[2]][47:40]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][47:40]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][47:40];
                    PSPIC[path_temp_d1[3]][47:40]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][47:40]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][47:40];
                    PSPIC[path_temp_d1[4]][47:40]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][47:40]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][47:40];
                    PSPIC[path_temp_d1[5]][47:40]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][47:40]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][47:40];
                    PSPIC[path_temp_d1[6]][47:40]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][47:40]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][47:40];
                    PSPIC[path_temp_d1[7]][47:40]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][47:40]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][47:40];
                    PSPIC[path_temp_d1[8]][47:40]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][47:40]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][47:40];
                    PSPIC[path_temp_d1[9]][47:40]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][47:40]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][47:40];
                    PSPIC[path_temp_d1[10]][47:40]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][47:40]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][47:40];
                    PSPIC[path_temp_d1[11]][47:40]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][47:40]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][47:40];
                    PSPIC[path_temp_d1[12]][47:40]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][47:40]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][47:40];
                    PSPIC[path_temp_d1[13]][47:40]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][47:40]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][47:40];
                    PSPIC[path_temp_d1[14]][47:40]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][47:40]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][47:40];
                    PSPIC[path_temp_d1[15]][47:40]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][47:40]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][47:40];
                    PSPIC[path_temp_d1[16]][47:40]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][47:40]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][47:40];
                    PSPIC[path_temp_d1[17]][47:40]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][47:40]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][47:40];
                    PSPIC[path_temp_d1[18]][47:40]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][47:40]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][47:40];
                    PSPIC[path_temp_d1[19]][47:40]<=(19==branching_pointer_old)?(PSPIC[path_temp_d1[19]][47:40]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][47:40];
                    PSPIC[path_temp_d1[20]][47:40]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][47:40]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][47:40];
                    PSPIC[path_temp_d1[21]][47:40]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][47:40]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][47:40];
                    PSPIC[path_temp_d1[22]][47:40]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][47:40]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][47:40];
                    PSPIC[path_temp_d1[23]][47:40]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][47:40]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][47:40];
                     end
                5'd6 : begin
                    PSPIC[path_temp_d1[0]][55:48]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][55:48]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][55:48];
                    PSPIC[path_temp_d1[1]][55:48]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][55:48]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][55:48];
                    PSPIC[path_temp_d1[2]][55:48]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][55:48]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][55:48];
                    PSPIC[path_temp_d1[3]][55:48]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][55:48]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][55:48];
                    PSPIC[path_temp_d1[4]][55:48]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][55:48]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][55:48];
                    PSPIC[path_temp_d1[5]][55:48]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][55:48]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][55:48];
                    PSPIC[path_temp_d1[6]][55:48]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][55:48]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][55:48];
                    PSPIC[path_temp_d1[7]][55:48]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][55:48]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][55:48];
                    PSPIC[path_temp_d1[8]][55:48]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][55:48]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][55:48];
                    PSPIC[path_temp_d1[9]][55:48]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][55:48]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][55:48];
                    PSPIC[path_temp_d1[10]][55:48]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][55:48]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][55:48];
                    PSPIC[path_temp_d1[11]][55:48]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][55:48]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][55:48];
                    PSPIC[path_temp_d1[12]][55:48]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][55:48]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][55:48];
                    PSPIC[path_temp_d1[13]][55:48]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][55:48]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][55:48];
                    PSPIC[path_temp_d1[14]][55:48]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][55:48]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][55:48];
                    PSPIC[path_temp_d1[15]][55:48]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][55:48]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][55:48];
                    PSPIC[path_temp_d1[16]][55:48]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][55:48]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][55:48];
                    PSPIC[path_temp_d1[17]][55:48]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][55:48]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][55:48];
                    PSPIC[path_temp_d1[18]][55:48]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][55:48]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][55:48];
                    PSPIC[path_temp_d1[19]][55:48]<=(19==branching_pointer_old)?(PSPIC[path_temp_d1[19]][55:48]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][55:48];
                    PSPIC[path_temp_d1[20]][55:48]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][55:48]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][55:48];
                    PSPIC[path_temp_d1[21]][55:48]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][55:48]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][55:48];
                    PSPIC[path_temp_d1[22]][55:48]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][55:48]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][55:48];
                    PSPIC[path_temp_d1[23]][55:48]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][55:48]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][55:48];end
                5'd7 : begin
                    PSPIC[path_temp_d1[0]][63:56]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][63:56]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][63:56];
                    PSPIC[path_temp_d1[1]][63:56]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][63:56]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][63:56];
                    PSPIC[path_temp_d1[2]][63:56]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][63:56]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][63:56];
                    PSPIC[path_temp_d1[3]][63:56]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][63:56]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][63:56];
                    PSPIC[path_temp_d1[4]][63:56]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][63:56]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][63:56];
                    PSPIC[path_temp_d1[5]][63:56]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][63:56]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][63:56];
                    PSPIC[path_temp_d1[6]][63:56]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][63:56]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][63:56];
                    PSPIC[path_temp_d1[7]][63:56]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][63:56]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][63:56];
                    PSPIC[path_temp_d1[8]][63:56]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][63:56]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][63:56];
                    PSPIC[path_temp_d1[9]][63:56]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][63:56]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][63:56];
                    PSPIC[path_temp_d1[10]][63:56]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][63:56]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][63:56];
                    PSPIC[path_temp_d1[11]][63:56]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][63:56]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][63:56];
                    PSPIC[path_temp_d1[12]][63:56]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][63:56]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][63:56];
                    PSPIC[path_temp_d1[13]][63:56]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][63:56]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][63:56];
                    PSPIC[path_temp_d1[14]][63:56]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][63:56]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][63:56];
                    PSPIC[path_temp_d1[15]][63:56]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][63:56]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][63:56];
                    PSPIC[path_temp_d1[16]][63:56]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][63:56]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][63:56];
                    PSPIC[path_temp_d1[17]][63:56]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][63:56]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][63:56];
                    PSPIC[path_temp_d1[18]][63:56]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][63:56]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][63:56];
                    PSPIC[path_temp_d1[19]][63:56]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][63:56]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][63:56];
                    PSPIC[path_temp_d1[20]][63:56]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][63:56]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][63:56];
                    PSPIC[path_temp_d1[21]][63:56]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][63:56]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][63:56];
                    PSPIC[path_temp_d1[22]][63:56]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][63:56]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][63:56];
                    PSPIC[path_temp_d1[23]][63:56]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][63:56]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][63:56];
                   // PSPIC[path_temp_d1[24]][63:56]<=(24>=branching_pointer_old)?(PSPIC[path_temp_d1[24]][63:56]+ps_invc_temp[24]):PSPIC[path_temp_d1[24]][63:56];
                     end
                5'd8 : begin
                    PSPIC[path_temp_d1[0]][71:64]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][71:64]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][71:64];
                    PSPIC[path_temp_d1[1]][71:64]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][71:64]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][71:64];
                    PSPIC[path_temp_d1[2]][71:64]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][71:64]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][71:64];
                    PSPIC[path_temp_d1[3]][71:64]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][71:64]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][71:64];
                    PSPIC[path_temp_d1[4]][71:64]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][71:64]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][71:64];
                    PSPIC[path_temp_d1[5]][71:64]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][71:64]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][71:64];
                    PSPIC[path_temp_d1[6]][71:64]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][71:64]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][71:64];
                    PSPIC[path_temp_d1[7]][71:64]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][71:64]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][71:64];
                    PSPIC[path_temp_d1[8]][71:64]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][71:64]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][71:64];
                    PSPIC[path_temp_d1[9]][71:64]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][71:64]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][71:64];
                    PSPIC[path_temp_d1[10]][71:64]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][71:64]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][71:64];
                    PSPIC[path_temp_d1[11]][71:64]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][71:64]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][71:64];
                    PSPIC[path_temp_d1[12]][71:64]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][71:64]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][71:64];
                    PSPIC[path_temp_d1[13]][71:64]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][71:64]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][71:64];
                    PSPIC[path_temp_d1[14]][71:64]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][71:64]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][71:64];
                    PSPIC[path_temp_d1[15]][71:64]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][71:64]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][71:64];
                    PSPIC[path_temp_d1[16]][71:64]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][71:64]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][71:64];
                    PSPIC[path_temp_d1[17]][71:64]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][71:64]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][71:64];
                    PSPIC[path_temp_d1[18]][71:64]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][71:64]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][71:64];
                    PSPIC[path_temp_d1[19]][71:64]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][71:64]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][71:64];
                    PSPIC[path_temp_d1[20]][71:64]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][71:64]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][71:64];
                    PSPIC[path_temp_d1[21]][71:64]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][71:64]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][71:64];
                    PSPIC[path_temp_d1[22]][71:64]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][71:64]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][71:64];
                    PSPIC[path_temp_d1[23]][71:64]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][71:64]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][71:64];
                     end
                5'd9 : begin
                    PSPIC[path_temp_d1[0]][79:72]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][79:72]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][79:72];
                    PSPIC[path_temp_d1[1]][79:72]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][79:72]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][79:72];
                    PSPIC[path_temp_d1[2]][79:72]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][79:72]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][79:72];
                    PSPIC[path_temp_d1[3]][79:72]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][79:72]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][79:72];
                    PSPIC[path_temp_d1[4]][79:72]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][79:72]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][79:72];
                    PSPIC[path_temp_d1[5]][79:72]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][79:72]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][79:72];
                    PSPIC[path_temp_d1[6]][79:72]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][79:72]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][79:72];
                    PSPIC[path_temp_d1[7]][79:72]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][79:72]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][79:72];
                    PSPIC[path_temp_d1[8]][79:72]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][79:72]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][79:72];
                    PSPIC[path_temp_d1[9]][79:72]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][79:72]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][79:72];
                    PSPIC[path_temp_d1[10]][79:72]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][79:72]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][79:72];
                    PSPIC[path_temp_d1[11]][79:72]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][79:72]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][79:72];
                    PSPIC[path_temp_d1[12]][79:72]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][79:72]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][79:72];
                    PSPIC[path_temp_d1[13]][79:72]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][79:72]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][79:72];
                    PSPIC[path_temp_d1[14]][79:72]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][79:72]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][79:72];
                    PSPIC[path_temp_d1[15]][79:72]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][79:72]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][79:72];
                    PSPIC[path_temp_d1[16]][79:72]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][79:72]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][79:72];
                    PSPIC[path_temp_d1[17]][79:72]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][79:72]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][79:72];
                    PSPIC[path_temp_d1[18]][79:72]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][79:72]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][79:72];
                    PSPIC[path_temp_d1[19]][79:72]<=(19==branching_pointer_old)?(PSPIC[path_temp_d1[19]][79:72]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][79:72];
                    PSPIC[path_temp_d1[20]][79:72]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][79:72]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][79:72];
                    PSPIC[path_temp_d1[21]][79:72]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][79:72]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][79:72];
                    PSPIC[path_temp_d1[22]][79:72]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][79:72]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][79:72];
                    PSPIC[path_temp_d1[23]][79:72]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][79:72]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][79:72];
                     end
                5'd10 : begin
                    PSPIC[path_temp_d1[0]][87:80]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][87:80]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][87:80];
                    PSPIC[path_temp_d1[1]][87:80]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][87:80]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][87:80];
                    PSPIC[path_temp_d1[2]][87:80]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][87:80]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][87:80];
                    PSPIC[path_temp_d1[3]][87:80]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][87:80]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][87:80];
                    PSPIC[path_temp_d1[4]][87:80]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][87:80]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][87:80];
                    PSPIC[path_temp_d1[5]][87:80]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][87:80]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][87:80];
                    PSPIC[path_temp_d1[6]][87:80]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][87:80]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][87:80];
                    PSPIC[path_temp_d1[7]][87:80]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][87:80]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][87:80];
                    PSPIC[path_temp_d1[8]][87:80]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][87:80]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][87:80];
                    PSPIC[path_temp_d1[9]][87:80]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][87:80]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][87:80];
                    PSPIC[path_temp_d1[10]][87:80]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][87:80]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][87:80];
                    PSPIC[path_temp_d1[11]][87:80]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][87:80]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][87:80];
                    PSPIC[path_temp_d1[12]][87:80]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][87:80]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][87:80];
                    PSPIC[path_temp_d1[13]][87:80]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][87:80]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][87:80];
                    PSPIC[path_temp_d1[14]][87:80]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][87:80]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][87:80];
                    PSPIC[path_temp_d1[15]][87:80]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][87:80]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][87:80];
                    PSPIC[path_temp_d1[16]][87:80]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][87:80]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][87:80];
                    PSPIC[path_temp_d1[17]][87:80]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][87:80]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][87:80];
                    PSPIC[path_temp_d1[18]][87:80]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][87:80]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][87:80];
                    PSPIC[path_temp_d1[19]][87:80]<=(19==branching_pointer_old)?(PSPIC[path_temp_d1[19]][87:80]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][87:80];
                    PSPIC[path_temp_d1[20]][87:80]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][87:80]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][87:80];
                    PSPIC[path_temp_d1[21]][87:80]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][87:80]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][87:80];
                    PSPIC[path_temp_d1[22]][87:80]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][87:80]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][87:80];
                    PSPIC[path_temp_d1[23]][87:80]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][87:80]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][87:80];
                     end
               5'd11 : begin
                    PSPIC[path_temp_d1[0]][95:88]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][95:88]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][95:88];
                    PSPIC[path_temp_d1[1]][95:88]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][95:88]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][95:88];
                    PSPIC[path_temp_d1[2]][95:88]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][95:88]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][95:88];
                    PSPIC[path_temp_d1[3]][95:88]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][95:88]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][95:88];
                    PSPIC[path_temp_d1[4]][95:88]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][95:88]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][95:88];
                    PSPIC[path_temp_d1[5]][95:88]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][95:88]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][95:88];
                    PSPIC[path_temp_d1[6]][95:88]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][95:88]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][95:88];
                    PSPIC[path_temp_d1[7]][95:88]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][95:88]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][95:88];
                    PSPIC[path_temp_d1[8]][95:88]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][95:88]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][95:88];
                    PSPIC[path_temp_d1[9]][95:88]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][95:88]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][95:88];
                    PSPIC[path_temp_d1[10]][95:88]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][95:88]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][95:88];
                    PSPIC[path_temp_d1[11]][95:88]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][95:88]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][95:88];
                    PSPIC[path_temp_d1[12]][95:88]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][95:88]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][95:88];
                    PSPIC[path_temp_d1[13]][95:88]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][95:88]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][95:88];
                    PSPIC[path_temp_d1[14]][95:88]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][95:88]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][95:88];
                    PSPIC[path_temp_d1[15]][95:88]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][95:88]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][95:88];
                    PSPIC[path_temp_d1[16]][95:88]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][95:88]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][95:88];
                    PSPIC[path_temp_d1[17]][95:88]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][95:88]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][95:88];
                    PSPIC[path_temp_d1[18]][95:88]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][95:88]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][95:88];
                    PSPIC[path_temp_d1[19]][95:88]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][95:88]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][95:88];
                    PSPIC[path_temp_d1[20]][95:88]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][95:88]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][95:88];
                    PSPIC[path_temp_d1[21]][95:88]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][95:88]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][95:88];
                    PSPIC[path_temp_d1[22]][95:88]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][95:88]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][95:88];
                    PSPIC[path_temp_d1[23]][95:88]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][95:88]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][95:88];
                     end//v1-zcu104*/
                5'd12 : begin
                    PSPIC[path_temp_d1[0]][103:96]<=(0>branching_pointer_old)?(PSPIC[path_temp_d1[0]][103:96]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][103:96];
                    PSPIC[path_temp_d1[1]][103:96]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][103:96]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][103:96];
                    PSPIC[path_temp_d1[2]][103:96]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][103:96]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][103:96];
                    PSPIC[path_temp_d1[3]][103:96]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][103:96]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][103:96];
                    PSPIC[path_temp_d1[4]][103:96]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][103:96]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][103:96];
                    PSPIC[path_temp_d1[5]][103:96]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][103:96]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][103:96];
                    PSPIC[path_temp_d1[6]][103:96]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][103:96]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][103:96];
                    PSPIC[path_temp_d1[7]][103:96]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][103:96]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][103:96];
                    PSPIC[path_temp_d1[8]][103:96]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][103:96]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][103:96];
                    PSPIC[path_temp_d1[9]][103:96]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][103:96]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][103:96];
                    PSPIC[path_temp_d1[10]][103:96]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][103:96]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][103:96];
                    PSPIC[path_temp_d1[11]][103:96]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][103:96]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][103:96];
                    PSPIC[path_temp_d1[12]][103:96]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][103:96]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][103:96];
                    PSPIC[path_temp_d1[13]][103:96]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][103:96]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][103:96];
                    PSPIC[path_temp_d1[14]][103:96]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][103:96]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][103:96];
                    PSPIC[path_temp_d1[15]][103:96]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][103:96]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][103:96];
                    PSPIC[path_temp_d1[16]][103:96]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][103:96]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][103:96];
                    PSPIC[path_temp_d1[17]][103:96]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][103:96]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][103:96];
                    PSPIC[path_temp_d1[18]][103:96]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][103:96]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][103:96];
                    PSPIC[path_temp_d1[19]][103:96]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][103:96]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][103:96];
                    PSPIC[path_temp_d1[20]][103:96]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][103:96]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][103:96];
                    PSPIC[path_temp_d1[21]][103:96]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][103:96]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][103:96];
                    PSPIC[path_temp_d1[22]][103:96]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][103:96]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][103:96];
                    PSPIC[path_temp_d1[23]][103:96]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][103:96]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][103:96];
                     end
                5'd13 : begin
                    PSPIC[path_temp_d1[0]][111:104]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][111:104]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][111:104];
                    PSPIC[path_temp_d1[1]][111:104]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][111:104]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][111:104];
                    PSPIC[path_temp_d1[2]][111:104]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][111:104]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][111:104];
                    PSPIC[path_temp_d1[3]][111:104]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][111:104]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][111:104];
                    PSPIC[path_temp_d1[4]][111:104]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][111:104]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][111:104];
                    PSPIC[path_temp_d1[5]][111:104]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][111:104]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][111:104];
                    PSPIC[path_temp_d1[6]][111:104]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][111:104]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][111:104];
                    PSPIC[path_temp_d1[7]][111:104]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][111:104]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][111:104];
                    PSPIC[path_temp_d1[8]][111:104]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][111:104]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][111:104];
                    PSPIC[path_temp_d1[9]][111:104]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][111:104]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][111:104];
                    PSPIC[path_temp_d1[10]][111:104]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][111:104]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][111:104];
                    PSPIC[path_temp_d1[11]][111:104]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][111:104]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][111:104];
                    PSPIC[path_temp_d1[12]][111:104]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][111:104]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][111:104];
                    PSPIC[path_temp_d1[13]][111:104]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][111:104]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][111:104];
                    PSPIC[path_temp_d1[14]][111:104]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][111:104]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][111:104];
                    PSPIC[path_temp_d1[15]][111:104]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][111:104]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][111:104];
                    PSPIC[path_temp_d1[16]][111:104]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][111:104]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][111:104];
                    PSPIC[path_temp_d1[17]][111:104]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][111:104]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][111:104];
                    PSPIC[path_temp_d1[18]][111:104]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][111:104]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][111:104];
                    PSPIC[path_temp_d1[19]][111:104]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][111:104]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][111:104];
  PSPIC[path_temp_d1[20]][111:104]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][111:104]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][111:104];
                    PSPIC[path_temp_d1[21]][111:104]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][111:104]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][111:104];
                    PSPIC[path_temp_d1[22]][111:104]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][111:104]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][111:104];
                    PSPIC[path_temp_d1[23]][111:104]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][111:104]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][111:104];end
                5'd14 : begin
                    PSPIC[path_temp_d1[0]][119:112]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][119:112]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][119:112];
                    PSPIC[path_temp_d1[1]][119:112]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][119:112]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][119:112];
                    PSPIC[path_temp_d1[2]][119:112]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][119:112]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][119:112];
                    PSPIC[path_temp_d1[3]][119:112]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][119:112]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][119:112];
                    PSPIC[path_temp_d1[4]][119:112]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][119:112]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][119:112];
                    PSPIC[path_temp_d1[5]][119:112]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][119:112]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][119:112];
                    PSPIC[path_temp_d1[6]][119:112]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][119:112]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][119:112];
                    PSPIC[path_temp_d1[7]][119:112]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][119:112]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][119:112];
                    PSPIC[path_temp_d1[8]][119:112]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][119:112]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][119:112];
                    PSPIC[path_temp_d1[9]][119:112]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][119:112]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][119:112];
                    PSPIC[path_temp_d1[10]][119:112]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][119:112]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][119:112];
                    PSPIC[path_temp_d1[11]][119:112]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][119:112]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][119:112];
                    PSPIC[path_temp_d1[12]][119:112]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][119:112]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][119:112];
                    PSPIC[path_temp_d1[13]][119:112]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][119:112]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][119:112];
                    PSPIC[path_temp_d1[14]][119:112]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][119:112]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][119:112];
                    PSPIC[path_temp_d1[15]][119:112]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][119:112]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][119:112];
                    PSPIC[path_temp_d1[16]][119:112]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][119:112]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][119:112];
                    PSPIC[path_temp_d1[17]][119:112]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][119:112]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][119:112];
                    PSPIC[path_temp_d1[18]][119:112]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][119:112]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][119:112];
                    PSPIC[path_temp_d1[19]][119:112]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][119:112]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][119:112];
                  PSPIC[path_temp_d1[20]][119:112]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][119:112]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][119:112];
                    PSPIC[path_temp_d1[21]][119:112]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][119:112]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][119:112];
                    PSPIC[path_temp_d1[22]][119:112]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][119:112]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][119:112];
                    PSPIC[path_temp_d1[23]][119:112]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][119:112]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][119:112];    end
               5'd15 : begin
                    PSPIC[path_temp_d1[0]][127:120]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][127:120]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][127:120];
                    PSPIC[path_temp_d1[1]][127:120]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][127:120]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][127:120];
                    PSPIC[path_temp_d1[2]][127:120]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][127:120]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][127:120];
                    PSPIC[path_temp_d1[3]][127:120]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][127:120]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][127:120];
                    PSPIC[path_temp_d1[4]][127:120]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][127:120]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][127:120];
                    PSPIC[path_temp_d1[5]][127:120]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][127:120]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][127:120];
                    PSPIC[path_temp_d1[6]][127:120]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][127:120]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][127:120];
                    PSPIC[path_temp_d1[7]][127:120]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][127:120]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][127:120];
                    PSPIC[path_temp_d1[8]][127:120]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][127:120]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][127:120];
                    PSPIC[path_temp_d1[9]][127:120]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][127:120]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][127:120];
                    PSPIC[path_temp_d1[10]][127:120]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][127:120]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][127:120];
                    PSPIC[path_temp_d1[11]][127:120]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][127:120]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][127:120];
                    PSPIC[path_temp_d1[12]][127:120]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][127:120]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][127:120];
                    PSPIC[path_temp_d1[13]][127:120]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][127:120]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][127:120];
                    PSPIC[path_temp_d1[14]][127:120]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][127:120]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][127:120];
                    PSPIC[path_temp_d1[15]][127:120]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][127:120]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][127:120];
                    PSPIC[path_temp_d1[16]][127:120]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][127:120]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][127:120];
                    PSPIC[path_temp_d1[17]][127:120]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][127:120]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][127:120];
                    PSPIC[path_temp_d1[18]][127:120]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][127:120]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][127:120];
                    PSPIC[path_temp_d1[19]][127:120]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][127:120]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][127:120];
 PSPIC[path_temp_d1[20]][127:120]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][127:120]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][127:120];
                    PSPIC[path_temp_d1[21]][127:120]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][127:120]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][127:120];
                    PSPIC[path_temp_d1[22]][127:120]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][127:120]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][127:120];
                    PSPIC[path_temp_d1[23]][127:120]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][127:120]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][127:120];
                     end
                5'd16 : begin
                    PSPIC[path_temp_d1[0]][135:128]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][135:128]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][135:128];
                    PSPIC[path_temp_d1[1]][135:128]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][135:128]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][135:128];
                    PSPIC[path_temp_d1[2]][135:128]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][135:128]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][135:128];
                    PSPIC[path_temp_d1[3]][135:128]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][135:128]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][135:128];
                    PSPIC[path_temp_d1[4]][135:128]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][135:128]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][135:128];
                    PSPIC[path_temp_d1[5]][135:128]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][135:128]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][135:128];
                    PSPIC[path_temp_d1[6]][135:128]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][135:128]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][135:128];
                    PSPIC[path_temp_d1[7]][135:128]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][135:128]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][135:128];
                    PSPIC[path_temp_d1[8]][135:128]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][135:128]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][135:128];
                    PSPIC[path_temp_d1[9]][135:128]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][135:128]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][135:128];
                    PSPIC[path_temp_d1[10]][135:128]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][135:128]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][135:128];
                    PSPIC[path_temp_d1[11]][135:128]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][135:128]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][135:128];
                    PSPIC[path_temp_d1[12]][135:128]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][135:128]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][135:128];
                    PSPIC[path_temp_d1[13]][135:128]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][135:128]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][135:128];
                    PSPIC[path_temp_d1[14]][135:128]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][135:128]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][135:128];
                    PSPIC[path_temp_d1[15]][135:128]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][135:128]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][135:128];
                    PSPIC[path_temp_d1[16]][135:128]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][135:128]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][135:128];
                    PSPIC[path_temp_d1[17]][135:128]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][135:128]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][135:128];
                    PSPIC[path_temp_d1[18]][135:128]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][135:128]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][135:128];
                    PSPIC[path_temp_d1[19]][135:128]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][135:128]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][135:128];
PSPIC[path_temp_d1[20]][135:128]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][135:128]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][135:128];
                    PSPIC[path_temp_d1[21]][135:128]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][135:128]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][135:128];
                    PSPIC[path_temp_d1[22]][135:128]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][135:128]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][135:128];
                    PSPIC[path_temp_d1[23]][135:128]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][135:128]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][135:128];
                     end
                5'd17 : begin
                    PSPIC[path_temp_d1[0]][143:136]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][143:136]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][143:136];
                    PSPIC[path_temp_d1[1]][143:136]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][143:136]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][143:136];
                    PSPIC[path_temp_d1[2]][143:136]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][143:136]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][143:136];
                    PSPIC[path_temp_d1[3]][143:136]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][143:136]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][143:136];
                    PSPIC[path_temp_d1[4]][143:136]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][143:136]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][143:136];
                    PSPIC[path_temp_d1[5]][143:136]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][143:136]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][143:136];
                    PSPIC[path_temp_d1[6]][143:136]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][143:136]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][143:136];
                    PSPIC[path_temp_d1[7]][143:136]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][143:136]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][143:136];
                    PSPIC[path_temp_d1[8]][143:136]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][143:136]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][143:136];
                    PSPIC[path_temp_d1[9]][143:136]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][143:136]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][143:136];
                    PSPIC[path_temp_d1[10]][143:136]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][143:136]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][143:136];
                    PSPIC[path_temp_d1[11]][143:136]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][143:136]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][143:136];
                    PSPIC[path_temp_d1[12]][143:136]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][143:136]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][143:136];
                    PSPIC[path_temp_d1[13]][143:136]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][143:136]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][143:136];
                    PSPIC[path_temp_d1[14]][143:136]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][143:136]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][143:136];
                    PSPIC[path_temp_d1[15]][143:136]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][143:136]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][143:136];
                    PSPIC[path_temp_d1[16]][143:136]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][143:136]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][143:136];
                    PSPIC[path_temp_d1[17]][143:136]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][143:136]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][143:136];
                    PSPIC[path_temp_d1[18]][143:136]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][143:136]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][143:136];
                    PSPIC[path_temp_d1[19]][143:136]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][143:136]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][143:136];
PSPIC[path_temp_d1[20]][143:136]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][143:136]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][143:136];
                    PSPIC[path_temp_d1[21]][143:136]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][143:136]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][143:136];
                    PSPIC[path_temp_d1[22]][143:136]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][143:136]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][143:136];
                    PSPIC[path_temp_d1[23]][143:136]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][143:136]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][143:136];
                     end
               5'd18 : begin
                    PSPIC[path_temp_d1[0]][151:144]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][151:144]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][151:144];
                    PSPIC[path_temp_d1[1]][151:144]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][151:144]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][151:144];
                    PSPIC[path_temp_d1[2]][151:144]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][151:144]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][151:144];
                    PSPIC[path_temp_d1[3]][151:144]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][151:144]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][151:144];
                    PSPIC[path_temp_d1[4]][151:144]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][151:144]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][151:144];
                    PSPIC[path_temp_d1[5]][151:144]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][151:144]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][151:144];
                    PSPIC[path_temp_d1[6]][151:144]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][151:144]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][151:144];
                    PSPIC[path_temp_d1[7]][151:144]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][151:144]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][151:144];
                    PSPIC[path_temp_d1[8]][151:144]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][151:144]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][151:144];
                    PSPIC[path_temp_d1[9]][151:144]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][151:144]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][151:144];
                    PSPIC[path_temp_d1[10]][151:144]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][151:144]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][151:144];
                    PSPIC[path_temp_d1[11]][151:144]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][151:144]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][151:144];
                    PSPIC[path_temp_d1[12]][151:144]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][151:144]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][151:144];
                    PSPIC[path_temp_d1[13]][151:144]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][151:144]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][151:144];
                    PSPIC[path_temp_d1[14]][151:144]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][151:144]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][151:144];
                    PSPIC[path_temp_d1[15]][151:144]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][151:144]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][151:144];
                    PSPIC[path_temp_d1[16]][151:144]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][151:144]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][151:144];
                    PSPIC[path_temp_d1[17]][151:144]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][151:144]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][151:144];
                    PSPIC[path_temp_d1[18]][151:144]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][151:144]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][151:144];
                    PSPIC[path_temp_d1[19]][151:144]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][151:144]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][151:144];
                    PSPIC[path_temp_d1[20]][151:144]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][151:144]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][151:144];
                    PSPIC[path_temp_d1[21]][151:144]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][151:144]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][151:144];
                    PSPIC[path_temp_d1[22]][151:144]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][151:144]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][151:144];
                    PSPIC[path_temp_d1[23]][151:144]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][151:144]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][151:144];
          end
                5'd19 : begin
                    PSPIC[path_temp_d1[0]][159:152]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][159:152]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][159:152];
                    PSPIC[path_temp_d1[1]][159:152]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][159:152]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][159:152];
                    PSPIC[path_temp_d1[2]][159:152]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][159:152]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][159:152];
                    PSPIC[path_temp_d1[3]][159:152]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][159:152]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][159:152];
                    PSPIC[path_temp_d1[4]][159:152]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][159:152]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][159:152];
                    PSPIC[path_temp_d1[5]][159:152]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][159:152]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][159:152];
                    PSPIC[path_temp_d1[6]][159:152]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][159:152]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][159:152];
                    PSPIC[path_temp_d1[7]][159:152]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][159:152]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][159:152];
                    PSPIC[path_temp_d1[8]][159:152]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][159:152]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][159:152];
                    PSPIC[path_temp_d1[9]][159:152]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][159:152]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][159:152];
                    PSPIC[path_temp_d1[10]][159:152]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][159:152]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][159:152];
                    PSPIC[path_temp_d1[11]][159:152]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][159:152]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][159:152];
                    PSPIC[path_temp_d1[12]][159:152]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][159:152]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][159:152];
                    PSPIC[path_temp_d1[13]][159:152]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][159:152]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][159:152];
                    PSPIC[path_temp_d1[14]][159:152]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][159:152]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][159:152];
                    PSPIC[path_temp_d1[15]][159:152]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][159:152]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][159:152];
                    PSPIC[path_temp_d1[16]][159:152]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][159:152]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][159:152];
                    PSPIC[path_temp_d1[17]][159:152]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][159:152]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][159:152];
                    PSPIC[path_temp_d1[18]][159:152]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][159:152]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][159:152];
                    PSPIC[path_temp_d1[19]][159:152]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][159:152]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][159:152];
                    PSPIC[path_temp_d1[20]][159:152]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][159:152]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][159:152];
                    PSPIC[path_temp_d1[21]][159:152]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][159:152]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][159:152];
                    PSPIC[path_temp_d1[22]][159:152]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][159:152]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][159:152];
                    PSPIC[path_temp_d1[23]][159:152]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][159:152]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][159:152];
       end
                5'd20 : begin
                    PSPIC[path_temp_d1[0]][167:160]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][167:160]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][167:160];
                    PSPIC[path_temp_d1[1]][167:160]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][167:160]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][167:160];
                    PSPIC[path_temp_d1[2]][167:160]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][167:160]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][167:160];
                    PSPIC[path_temp_d1[3]][167:160]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][167:160]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][167:160];
                    PSPIC[path_temp_d1[4]][167:160]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][167:160]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][167:160];
                    PSPIC[path_temp_d1[5]][167:160]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][167:160]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][167:160];
                    PSPIC[path_temp_d1[6]][167:160]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][167:160]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][167:160];
                    PSPIC[path_temp_d1[7]][167:160]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][167:160]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][167:160];
                    PSPIC[path_temp_d1[8]][167:160]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][167:160]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][167:160];
                    PSPIC[path_temp_d1[9]][167:160]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][167:160]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][167:160];
                    PSPIC[path_temp_d1[10]][167:160]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][167:160]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][167:160];
                    PSPIC[path_temp_d1[11]][167:160]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][167:160]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][167:160];
                    PSPIC[path_temp_d1[12]][167:160]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][167:160]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][167:160];
                    PSPIC[path_temp_d1[13]][167:160]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][167:160]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][167:160];
                    PSPIC[path_temp_d1[14]][167:160]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][167:160]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][167:160];
                    PSPIC[path_temp_d1[15]][167:160]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][167:160]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][167:160];
                    PSPIC[path_temp_d1[16]][167:160]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][167:160]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][167:160];
                    PSPIC[path_temp_d1[17]][167:160]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][167:160]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][167:160];
                    PSPIC[path_temp_d1[18]][167:160]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][167:160]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][167:160];
                    PSPIC[path_temp_d1[19]][167:160]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][167:160]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][167:160];
                    PSPIC[path_temp_d1[20]][167:160]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][167:160]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][167:160];
                    PSPIC[path_temp_d1[21]][167:160]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][167:160]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][167:160];
                    PSPIC[path_temp_d1[22]][167:160]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][167:160]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][167:160];
                    PSPIC[path_temp_d1[23]][167:160]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][167:160]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][167:160];
   end
                5'd21 : begin
                    PSPIC[path_temp_d1[0]][175:168]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][175:168]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][175:168];
                    PSPIC[path_temp_d1[1]][175:168]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][175:168]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][175:168];
                    PSPIC[path_temp_d1[2]][175:168]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][175:168]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][175:168];
                    PSPIC[path_temp_d1[3]][175:168]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][175:168]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][175:168];
                    PSPIC[path_temp_d1[4]][175:168]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][175:168]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][175:168];
                    PSPIC[path_temp_d1[5]][175:168]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][175:168]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][175:168];
                    PSPIC[path_temp_d1[6]][175:168]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][175:168]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][175:168];
                    PSPIC[path_temp_d1[7]][175:168]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][175:168]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][175:168];
                    PSPIC[path_temp_d1[8]][175:168]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][175:168]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][175:168];
                    PSPIC[path_temp_d1[9]][175:168]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][175:168]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][175:168];
                    PSPIC[path_temp_d1[10]][175:168]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][175:168]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][175:168];
                    PSPIC[path_temp_d1[11]][175:168]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][175:168]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][175:168];
                    PSPIC[path_temp_d1[12]][175:168]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][175:168]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][175:168];
                    PSPIC[path_temp_d1[13]][175:168]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][175:168]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][175:168];
                    PSPIC[path_temp_d1[14]][175:168]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][175:168]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][175:168];
                    PSPIC[path_temp_d1[15]][175:168]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][175:168]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][175:168];
                    PSPIC[path_temp_d1[16]][175:168]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][175:168]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][175:168];
                    PSPIC[path_temp_d1[17]][175:168]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][175:168]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][175:168];
                    PSPIC[path_temp_d1[18]][175:168]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][175:168]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][175:168];
                    PSPIC[path_temp_d1[19]][175:168]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][175:168]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][175:168];
                    PSPIC[path_temp_d1[20]][175:168]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][175:168]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][175:168];
                    PSPIC[path_temp_d1[21]][175:168]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][175:168]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][175:168];
                    PSPIC[path_temp_d1[22]][175:168]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][175:168]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][175:168];
                    PSPIC[path_temp_d1[23]][175:168]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][175:168]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][175:168];
 end
                5'd22 : begin
                    PSPIC[path_temp_d1[0]][183:176]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][183:176]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][183:176];
                    PSPIC[path_temp_d1[1]][183:176]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][183:176]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][183:176];
                    PSPIC[path_temp_d1[2]][183:176]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][183:176]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][183:176];
                    PSPIC[path_temp_d1[3]][183:176]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][183:176]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][183:176];
                    PSPIC[path_temp_d1[4]][183:176]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][183:176]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][183:176];
                    PSPIC[path_temp_d1[5]][183:176]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][183:176]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][183:176];
                    PSPIC[path_temp_d1[6]][183:176]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][183:176]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][183:176];
                    PSPIC[path_temp_d1[7]][183:176]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][183:176]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][183:176];
                    PSPIC[path_temp_d1[8]][183:176]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][183:176]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][183:176];
                    PSPIC[path_temp_d1[9]][183:176]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][183:176]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][183:176];
                    PSPIC[path_temp_d1[10]][183:176]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][183:176]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][183:176];
                    PSPIC[path_temp_d1[11]][183:176]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][183:176]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][183:176];
                    PSPIC[path_temp_d1[12]][183:176]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][183:176]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][183:176];
                    PSPIC[path_temp_d1[13]][183:176]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][183:176]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][183:176];
                    PSPIC[path_temp_d1[14]][183:176]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][183:176]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][183:176];
                    PSPIC[path_temp_d1[15]][183:176]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][183:176]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][183:176];
                    PSPIC[path_temp_d1[16]][183:176]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][183:176]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][183:176];
                    PSPIC[path_temp_d1[17]][183:176]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][183:176]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][183:176];
                    PSPIC[path_temp_d1[18]][183:176]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][183:176]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][183:176];
                    PSPIC[path_temp_d1[19]][183:176]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][183:176]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][183:176];
                    PSPIC[path_temp_d1[20]][183:176]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][183:176]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][183:176];
                    PSPIC[path_temp_d1[21]][183:176]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][183:176]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][183:176];
                    PSPIC[path_temp_d1[22]][183:176]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][183:176]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][183:176];
                    PSPIC[path_temp_d1[23]][183:176]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][183:176]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][183:176];
                      end
                5'd23 : begin
                    PSPIC[path_temp_d1[0]][191:184]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][191:184]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][191:184];
                    PSPIC[path_temp_d1[1]][191:184]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][191:184]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][191:184];
                    PSPIC[path_temp_d1[2]][191:184]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][191:184]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][191:184];
                    PSPIC[path_temp_d1[3]][191:184]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][191:184]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][191:184];
                    PSPIC[path_temp_d1[4]][191:184]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][191:184]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][191:184];
                    PSPIC[path_temp_d1[5]][191:184]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][191:184]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][191:184];
                    PSPIC[path_temp_d1[6]][191:184]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][191:184]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][191:184];
                    PSPIC[path_temp_d1[7]][191:184]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][191:184]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][191:184];
                    PSPIC[path_temp_d1[8]][191:184]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][191:184]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][191:184];
                    PSPIC[path_temp_d1[9]][191:184]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][191:184]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][191:184];
                    PSPIC[path_temp_d1[10]][191:184]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][191:184]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][191:184];
                    PSPIC[path_temp_d1[11]][191:184]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][191:184]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][191:184];
                    PSPIC[path_temp_d1[12]][191:184]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][191:184]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][191:184];
                    PSPIC[path_temp_d1[13]][191:184]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][191:184]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][191:184];
                    PSPIC[path_temp_d1[14]][191:184]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][191:184]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][191:184];
                    PSPIC[path_temp_d1[15]][191:184]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][191:184]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][191:184];
                    PSPIC[path_temp_d1[16]][191:184]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][191:184]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][191:184];
                    PSPIC[path_temp_d1[17]][191:184]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][191:184]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][191:184];
                    PSPIC[path_temp_d1[18]][191:184]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][191:184]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][191:184];
                    PSPIC[path_temp_d1[19]][191:184]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][191:184]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][191:184];
                    PSPIC[path_temp_d1[20]][191:184]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][191:184]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][191:184];
                    PSPIC[path_temp_d1[21]][191:184]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][191:184]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][191:184];
                    PSPIC[path_temp_d1[22]][191:184]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][191:184]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][191:184];
                    PSPIC[path_temp_d1[23]][191:184]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][191:184]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][191:184];
                     end
                5'd24 : begin
                    PSPIC[path_temp_d1[0]][199:192]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][199:192]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][199:192];
                    PSPIC[path_temp_d1[1]][199:192]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][199:192]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][199:192];
                    PSPIC[path_temp_d1[2]][199:192]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][199:192]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][199:192];
                    PSPIC[path_temp_d1[3]][199:192]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][199:192]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][199:192];
                    PSPIC[path_temp_d1[4]][199:192]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][199:192]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][199:192];
                    PSPIC[path_temp_d1[5]][199:192]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][199:192]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][199:192];
                    PSPIC[path_temp_d1[6]][199:192]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][199:192]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][199:192];
                    PSPIC[path_temp_d1[7]][199:192]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][199:192]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][199:192];
                    PSPIC[path_temp_d1[8]][199:192]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][199:192]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][199:192];
                    PSPIC[path_temp_d1[9]][199:192]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][199:192]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][199:192];
                    PSPIC[path_temp_d1[10]][199:192]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][199:192]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][199:192];
                    PSPIC[path_temp_d1[11]][199:192]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][199:192]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][199:192];
                    PSPIC[path_temp_d1[12]][199:192]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][199:192]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][199:192];
                    PSPIC[path_temp_d1[13]][199:192]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][199:192]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][199:192];
                    PSPIC[path_temp_d1[14]][199:192]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][199:192]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][199:192];
                    PSPIC[path_temp_d1[15]][199:192]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][199:192]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][199:192];
                    PSPIC[path_temp_d1[16]][199:192]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][199:192]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][199:192];
                    PSPIC[path_temp_d1[17]][199:192]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][199:192]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][199:192];
                    PSPIC[path_temp_d1[18]][199:192]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][199:192]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][199:192];
                    PSPIC[path_temp_d1[19]][199:192]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][199:192]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][199:192];
                    PSPIC[path_temp_d1[20]][199:192]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][199:192]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][199:192];
                    PSPIC[path_temp_d1[21]][199:192]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][199:192]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][199:192];
                    PSPIC[path_temp_d1[22]][199:192]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][199:192]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][199:192];
                    PSPIC[path_temp_d1[23]][199:192]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][199:192]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][199:192];
                     end
               5'd25 : begin
                    PSPIC[path_temp_d1[0]][207:200]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][207:200]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][207:200];
                    PSPIC[path_temp_d1[1]][207:200]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][207:200]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][207:200];
                    PSPIC[path_temp_d1[2]][207:200]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][207:200]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][207:200];
                    PSPIC[path_temp_d1[3]][207:200]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][207:200]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][207:200];
                    PSPIC[path_temp_d1[4]][207:200]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][207:200]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][207:200];
                    PSPIC[path_temp_d1[5]][207:200]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][207:200]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][207:200];
                    PSPIC[path_temp_d1[6]][207:200]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][207:200]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][207:200];
                    PSPIC[path_temp_d1[7]][207:200]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][207:200]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][207:200];
                    PSPIC[path_temp_d1[8]][207:200]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][207:200]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][207:200];
                    PSPIC[path_temp_d1[9]][207:200]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][207:200]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][207:200];
                    PSPIC[path_temp_d1[10]][207:200]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][207:200]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][207:200];
                    PSPIC[path_temp_d1[11]][207:200]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][207:200]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][207:200];
                    PSPIC[path_temp_d1[12]][207:200]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][207:200]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][207:200];
                    PSPIC[path_temp_d1[13]][207:200]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][207:200]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][207:200];
                    PSPIC[path_temp_d1[14]][207:200]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][207:200]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][207:200];
                    PSPIC[path_temp_d1[15]][207:200]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][207:200]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][207:200];
                    PSPIC[path_temp_d1[16]][207:200]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][207:200]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][207:200];
                    PSPIC[path_temp_d1[17]][207:200]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][207:200]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][207:200];
                    PSPIC[path_temp_d1[18]][207:200]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][207:200]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][207:200];
                    PSPIC[path_temp_d1[19]][207:200]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][207:200]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][207:200];
                    PSPIC[path_temp_d1[20]][207:200]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][207:200]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][207:200];
                    PSPIC[path_temp_d1[21]][207:200]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][207:200]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][207:200];
                    PSPIC[path_temp_d1[22]][207:200]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][207:200]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][207:200];
                    PSPIC[path_temp_d1[23]][207:200]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][207:200]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][207:200];
                     end
                5'd26 : begin
                    PSPIC[path_temp_d1[0]][215:208]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][215:208]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][215:208];
                    PSPIC[path_temp_d1[1]][215:208]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][215:208]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][215:208];
                    PSPIC[path_temp_d1[2]][215:208]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][215:208]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][215:208];
                    PSPIC[path_temp_d1[3]][215:208]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][215:208]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][215:208];
                    PSPIC[path_temp_d1[4]][215:208]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][215:208]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][215:208];
                    PSPIC[path_temp_d1[5]][215:208]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][215:208]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][215:208];
                    PSPIC[path_temp_d1[6]][215:208]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][215:208]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][215:208];
                    PSPIC[path_temp_d1[7]][215:208]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][215:208]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][215:208];
                    PSPIC[path_temp_d1[8]][215:208]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][215:208]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][215:208];
                    PSPIC[path_temp_d1[9]][215:208]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][215:208]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][215:208];
                    PSPIC[path_temp_d1[10]][215:208]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][215:208]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][215:208];
                    PSPIC[path_temp_d1[11]][215:208]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][215:208]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][215:208];
                    PSPIC[path_temp_d1[12]][215:208]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][215:208]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][215:208];
                    PSPIC[path_temp_d1[13]][215:208]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][215:208]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][215:208];
                    PSPIC[path_temp_d1[14]][215:208]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][215:208]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][215:208];
                    PSPIC[path_temp_d1[15]][215:208]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][215:208]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][215:208];
                    PSPIC[path_temp_d1[16]][215:208]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][215:208]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][215:208];
                    PSPIC[path_temp_d1[17]][215:208]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][215:208]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][215:208];
                    PSPIC[path_temp_d1[18]][215:208]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][215:208]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][215:208];
                    PSPIC[path_temp_d1[19]][215:208]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][215:208]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][215:208];
                    PSPIC[path_temp_d1[20]][215:208]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][215:208]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][215:208];
                    PSPIC[path_temp_d1[21]][215:208]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][215:208]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][215:208];
                    PSPIC[path_temp_d1[22]][215:208]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][215:208]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][215:208];
                    PSPIC[path_temp_d1[23]][215:208]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][215:208]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][215:208];
                     end
                5'd27 : begin
                    PSPIC[path_temp_d1[0]][223:216]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][223:216]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][223:216];
                    PSPIC[path_temp_d1[1]][223:216]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][223:216]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][223:216];
                    PSPIC[path_temp_d1[2]][223:216]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][223:216]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][223:216];
                    PSPIC[path_temp_d1[3]][223:216]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][223:216]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][223:216];
                    PSPIC[path_temp_d1[4]][223:216]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][223:216]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][223:216];
                    PSPIC[path_temp_d1[5]][223:216]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][223:216]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][223:216];
                    PSPIC[path_temp_d1[6]][223:216]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][223:216]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][223:216];
                    PSPIC[path_temp_d1[7]][223:216]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][223:216]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][223:216];
                    PSPIC[path_temp_d1[8]][223:216]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][223:216]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][223:216];
                    PSPIC[path_temp_d1[9]][223:216]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][223:216]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][223:216];
                    PSPIC[path_temp_d1[10]][223:216]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][223:216]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][223:216];
                    PSPIC[path_temp_d1[11]][223:216]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][223:216]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][223:216];
                    PSPIC[path_temp_d1[12]][223:216]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][223:216]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][223:216];
                    PSPIC[path_temp_d1[13]][223:216]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][223:216]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][223:216];
                    PSPIC[path_temp_d1[14]][223:216]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][223:216]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][223:216];
                    PSPIC[path_temp_d1[15]][223:216]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][223:216]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][223:216];
                    PSPIC[path_temp_d1[16]][223:216]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][223:216]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][223:216];
                    PSPIC[path_temp_d1[17]][223:216]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][223:216]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][223:216];
                    PSPIC[path_temp_d1[18]][223:216]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][223:216]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][223:216];
                    PSPIC[path_temp_d1[19]][223:216]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][223:216]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][223:216];
                    PSPIC[path_temp_d1[20]][223:216]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][223:216]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][223:216];
                    PSPIC[path_temp_d1[21]][223:216]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][223:216]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][223:216];
                    PSPIC[path_temp_d1[22]][223:216]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][223:216]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][223:216];
                    PSPIC[path_temp_d1[23]][223:216]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][223:216]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][223:216];
                     end
                5'd28 : begin
                    PSPIC[path_temp_d1[0]][231:224]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][231:224]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][231:224];
                    PSPIC[path_temp_d1[1]][231:224]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][231:224]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][231:224];
                    PSPIC[path_temp_d1[2]][231:224]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][231:224]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][231:224];
                    PSPIC[path_temp_d1[3]][231:224]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][231:224]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][231:224];
                    PSPIC[path_temp_d1[4]][231:224]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][231:224]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][231:224];
                    PSPIC[path_temp_d1[5]][231:224]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][231:224]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][231:224];
                    PSPIC[path_temp_d1[6]][231:224]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][231:224]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][231:224];
                    PSPIC[path_temp_d1[7]][231:224]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][231:224]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][231:224];
                    PSPIC[path_temp_d1[8]][231:224]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][231:224]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][231:224];
                    PSPIC[path_temp_d1[9]][231:224]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][231:224]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][231:224];
                    PSPIC[path_temp_d1[10]][231:224]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][231:224]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][231:224];
                    PSPIC[path_temp_d1[11]][231:224]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][231:224]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][231:224];
                    PSPIC[path_temp_d1[12]][231:224]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][231:224]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][231:224];
                    PSPIC[path_temp_d1[13]][231:224]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][231:224]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][231:224];
                    PSPIC[path_temp_d1[14]][231:224]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][231:224]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][231:224];
                    PSPIC[path_temp_d1[15]][231:224]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][231:224]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][231:224];
                    PSPIC[path_temp_d1[16]][231:224]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][231:224]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][231:224];
                    PSPIC[path_temp_d1[17]][231:224]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][231:224]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][231:224];
                    PSPIC[path_temp_d1[18]][231:224]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][231:224]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][231:224];
                    PSPIC[path_temp_d1[19]][231:224]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][231:224]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][231:224];
                    PSPIC[path_temp_d1[20]][231:224]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][231:224]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][231:224];
                    PSPIC[path_temp_d1[21]][231:224]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][231:224]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][231:224];
                    PSPIC[path_temp_d1[22]][231:224]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][231:224]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][231:224];
                    PSPIC[path_temp_d1[23]][231:224]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][231:224]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][231:224];
                     end
                5'd29 : begin
                    PSPIC[path_temp_d1[0]][239:232]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][239:232]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][239:232];
                    PSPIC[path_temp_d1[1]][239:232]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][239:232]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][239:232];
                    PSPIC[path_temp_d1[2]][239:232]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][239:232]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][239:232];
                    PSPIC[path_temp_d1[3]][239:232]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][239:232]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][239:232];
                    PSPIC[path_temp_d1[4]][239:232]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][239:232]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][239:232];
                    PSPIC[path_temp_d1[5]][239:232]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][239:232]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][239:232];
                    PSPIC[path_temp_d1[6]][239:232]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][239:232]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][239:232];
                    PSPIC[path_temp_d1[7]][239:232]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][239:232]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][239:232];
                    PSPIC[path_temp_d1[8]][239:232]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][239:232]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][239:232];
                    PSPIC[path_temp_d1[9]][239:232]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][239:232]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][239:232];
                    PSPIC[path_temp_d1[10]][239:232]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][239:232]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][239:232];
                    PSPIC[path_temp_d1[11]][239:232]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][239:232]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][239:232];
                    PSPIC[path_temp_d1[12]][239:232]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][239:232]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][239:232];
                    PSPIC[path_temp_d1[13]][239:232]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][239:232]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][239:232];
                    PSPIC[path_temp_d1[14]][239:232]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][239:232]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][239:232];
                    PSPIC[path_temp_d1[15]][239:232]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][239:232]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][239:232];
                    PSPIC[path_temp_d1[16]][239:232]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][239:232]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][239:232];
                    PSPIC[path_temp_d1[17]][239:232]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][239:232]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][239:232];
                    PSPIC[path_temp_d1[18]][239:232]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][239:232]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][239:232];
                    PSPIC[path_temp_d1[19]][239:232]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][239:232]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][239:232];
                    PSPIC[path_temp_d1[20]][239:232]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][239:232]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][239:232];
                    PSPIC[path_temp_d1[21]][239:232]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][239:232]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][239:232];
                    PSPIC[path_temp_d1[22]][239:232]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][239:232]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][239:232];
                    PSPIC[path_temp_d1[23]][239:232]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][239:232]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][239:232];
                     end
                5'd30 : begin
                    PSPIC[path_temp_d1[0]][247:240]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][247:240]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][247:240];
                    PSPIC[path_temp_d1[1]][247:240]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][247:240]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][247:240];
                    PSPIC[path_temp_d1[2]][247:240]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][247:240]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][247:240];
                    PSPIC[path_temp_d1[3]][247:240]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][247:240]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][247:240];
                    PSPIC[path_temp_d1[4]][247:240]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][247:240]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][247:240];
                    PSPIC[path_temp_d1[5]][247:240]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][247:240]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][247:240];
                    PSPIC[path_temp_d1[6]][247:240]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][247:240]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][247:240];
                    PSPIC[path_temp_d1[7]][247:240]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][247:240]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][247:240];
                    PSPIC[path_temp_d1[8]][247:240]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][247:240]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][247:240];
                    PSPIC[path_temp_d1[9]][247:240]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][247:240]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][247:240];
                    PSPIC[path_temp_d1[10]][247:240]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][247:240]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][247:240];
                    PSPIC[path_temp_d1[11]][247:240]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][247:240]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][247:240];
                    PSPIC[path_temp_d1[12]][247:240]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][247:240]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][247:240];
                    PSPIC[path_temp_d1[13]][247:240]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][247:240]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][247:240];
                    PSPIC[path_temp_d1[14]][247:240]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][247:240]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][247:240];
                    PSPIC[path_temp_d1[15]][247:240]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][247:240]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][247:240];
                    PSPIC[path_temp_d1[16]][247:240]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][247:240]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][247:240];
                    PSPIC[path_temp_d1[17]][247:240]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][247:240]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][247:240];
                    PSPIC[path_temp_d1[18]][247:240]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][247:240]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][247:240];
                    PSPIC[path_temp_d1[19]][247:240]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][247:240]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][247:240];
                    PSPIC[path_temp_d1[20]][247:240]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][247:240]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][247:240];
                    PSPIC[path_temp_d1[21]][247:240]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][247:240]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][247:240];
                    PSPIC[path_temp_d1[22]][247:240]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][247:240]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][247:240];
                    PSPIC[path_temp_d1[23]][247:240]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][247:240]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][247:240];
                     end
                default : begin
                    PSPIC[path_temp_d1[0]][255:248]<=(0>=branching_pointer_old)?(PSPIC[path_temp_d1[0]][255:248]+ps_invc_temp[0]):PSPIC[path_temp_d1[0]][255:248];
                    PSPIC[path_temp_d1[1]][255:248]<=(1>=branching_pointer_old)?(PSPIC[path_temp_d1[1]][255:248]+ps_invc_temp[1]):PSPIC[path_temp_d1[1]][255:248];
                    PSPIC[path_temp_d1[2]][255:248]<=(2>=branching_pointer_old)?(PSPIC[path_temp_d1[2]][255:248]+ps_invc_temp[2]):PSPIC[path_temp_d1[2]][255:248];
                    PSPIC[path_temp_d1[3]][255:248]<=(3>=branching_pointer_old)?(PSPIC[path_temp_d1[3]][255:248]+ps_invc_temp[3]):PSPIC[path_temp_d1[3]][255:248];
                    PSPIC[path_temp_d1[4]][255:248]<=(4>=branching_pointer_old)?(PSPIC[path_temp_d1[4]][255:248]+ps_invc_temp[4]):PSPIC[path_temp_d1[4]][255:248];
                    PSPIC[path_temp_d1[5]][255:248]<=(5>=branching_pointer_old)?(PSPIC[path_temp_d1[5]][255:248]+ps_invc_temp[5]):PSPIC[path_temp_d1[5]][255:248];
                    PSPIC[path_temp_d1[6]][255:248]<=(6>=branching_pointer_old)?(PSPIC[path_temp_d1[6]][255:248]+ps_invc_temp[6]):PSPIC[path_temp_d1[6]][255:248];
                    PSPIC[path_temp_d1[7]][255:248]<=(7>=branching_pointer_old)?(PSPIC[path_temp_d1[7]][255:248]+ps_invc_temp[7]):PSPIC[path_temp_d1[7]][255:248];
                    PSPIC[path_temp_d1[8]][255:248]<=(8>=branching_pointer_old)?(PSPIC[path_temp_d1[8]][255:248]+ps_invc_temp[8]):PSPIC[path_temp_d1[8]][255:248];
                    PSPIC[path_temp_d1[9]][255:248]<=(9>=branching_pointer_old)?(PSPIC[path_temp_d1[9]][255:248]+ps_invc_temp[9]):PSPIC[path_temp_d1[9]][255:248];
                    PSPIC[path_temp_d1[10]][255:248]<=(10>=branching_pointer_old)?(PSPIC[path_temp_d1[10]][255:248]+ps_invc_temp[10]):PSPIC[path_temp_d1[10]][255:248];
                    PSPIC[path_temp_d1[11]][255:248]<=(11>=branching_pointer_old)?(PSPIC[path_temp_d1[11]][255:248]+ps_invc_temp[11]):PSPIC[path_temp_d1[11]][255:248];
                    PSPIC[path_temp_d1[12]][255:248]<=(12>=branching_pointer_old)?(PSPIC[path_temp_d1[12]][255:248]+ps_invc_temp[12]):PSPIC[path_temp_d1[12]][255:248];
                    PSPIC[path_temp_d1[13]][255:248]<=(13>=branching_pointer_old)?(PSPIC[path_temp_d1[13]][255:248]+ps_invc_temp[13]):PSPIC[path_temp_d1[13]][255:248];
                    PSPIC[path_temp_d1[14]][255:248]<=(14>=branching_pointer_old)?(PSPIC[path_temp_d1[14]][255:248]+ps_invc_temp[14]):PSPIC[path_temp_d1[14]][255:248];
                    PSPIC[path_temp_d1[15]][255:248]<=(15>=branching_pointer_old)?(PSPIC[path_temp_d1[15]][255:248]+ps_invc_temp[15]):PSPIC[path_temp_d1[15]][255:248];
                    PSPIC[path_temp_d1[16]][255:248]<=(16>=branching_pointer_old)?(PSPIC[path_temp_d1[16]][255:248]+ps_invc_temp[16]):PSPIC[path_temp_d1[16]][255:248];
                    PSPIC[path_temp_d1[17]][255:248]<=(17>=branching_pointer_old)?(PSPIC[path_temp_d1[17]][255:248]+ps_invc_temp[17]):PSPIC[path_temp_d1[17]][255:248];
                    PSPIC[path_temp_d1[18]][255:248]<=(18>=branching_pointer_old)?(PSPIC[path_temp_d1[18]][255:248]+ps_invc_temp[18]):PSPIC[path_temp_d1[18]][255:248];
                    PSPIC[path_temp_d1[19]][255:248]<=(19>=branching_pointer_old)?(PSPIC[path_temp_d1[19]][255:248]+ps_invc_temp[19]):PSPIC[path_temp_d1[19]][255:248];
                    PSPIC[path_temp_d1[20]][255:248]<=(20>=branching_pointer_old)?(PSPIC[path_temp_d1[20]][255:248]+ps_invc_temp[20]):PSPIC[path_temp_d1[20]][255:248];
                    PSPIC[path_temp_d1[21]][255:248]<=(21>=branching_pointer_old)?(PSPIC[path_temp_d1[21]][255:248]+ps_invc_temp[21]):PSPIC[path_temp_d1[21]][255:248];
                    PSPIC[path_temp_d1[22]][255:248]<=(22>=branching_pointer_old)?(PSPIC[path_temp_d1[22]][255:248]+ps_invc_temp[22]):PSPIC[path_temp_d1[22]][255:248];
                    PSPIC[path_temp_d1[23]][255:248]<=(23==branching_pointer_old)?(PSPIC[path_temp_d1[23]][255:248]+ps_invc_temp[23]):PSPIC[path_temp_d1[23]][255:248];

                    end




                endcase 				 			       
end
else;
end

hit_path hit_path_1(
  .clk(clk),
  .reset(reset),
  .write_en(hit_wr_en), //st7_d2
  .addr(path_addr_d1), // from match_addr - was taking addr of func 16-11-2020
  .data_out0(hit_out0),
  .data_out1(hit_out1),
  .data_out2(hit_out2),
  .data_out3(hit_out3),
  .data_out4(hit_out4),
  .data_out5(hit_out5),
  .data_out6(hit_out6),
  .data_out7(hit_out7),
  .data_out8(hit_out8),
  .data_out9(hit_out9),
  .data_out10(hit_out10),
  .data_out11(hit_out11),
  .data_out12(hit_out12),
  .data_out13(hit_out13),
  .data_out14(hit_out14),
  .data_out15(hit_out15),
  .data_out16(hit_out16),
  .data_out17(hit_out17),
  .data_out18(hit_out18),
  .data_out19(hit_out19),
  .data_out20(hit_out20),
  .data_out21(hit_out21),
  .data_out22(hit_out22),
  .data_out23(hit_out23),
  .data_out24(hit_out24),
  .data_out25(hit_out25),
  .data_out26(hit_out26),
  .data_out27(hit_out27),
  .data_out28(hit_out28),
  .data_out29(hit_out29),
  .data_out30(hit_out30),
  .data_out31(hit_out31)
	); 



assign pcam_out0 = cam[0];
assign pcam_out1 = cam[1];
assign pcam_out2 = cam[2];
assign pcam_out3 = cam[3];
assign pcam_out4 = cam[4];
assign pcam_out5 = cam[5];
assign pcam_out6 = cam[6];
assign pcam_out7 = cam[7];
assign pcam_out8 = cam[8];
assign pcam_out9 = cam[9];
assign pcam_out10 = cam[10];
assign pcam_out11 = cam[11];
assign pcam_out12 = cam[12];
assign pcam_out13 = cam[13];
assign pcam_out14 = cam[14];
assign pcam_out15 = cam[15];
assign pcam_out16 = cam[16];
assign pcam_out17 = cam[17];
assign pcam_out18 = cam[18];
assign pcam_out19 = cam[19];
assign pcam_out20 = cam[20];
assign pcam_out21 = cam[21];
assign pcam_out22 = cam[22];
assign pcam_out23 = cam[23];
assign pcam_out24 = cam[24];
assign pcam_out25 = cam[25];
assign pcam_out26 = cam[26];
assign pcam_out27 = cam[27];
assign pcam_out28 = cam[28];
assign pcam_out29 = cam[29];
assign pcam_out30 = cam[30];
assign pcam_out31 = cam[31];




assign PSPIC0 = { PSPIC[0][255:248], PSPIC[0][247:240], PSPIC[0][239:232], PSPIC[0][231:224], PSPIC[0][223:216], PSPIC[0][215:208], PSPIC[0][207:200], PSPIC[0][199:192], PSPIC[0][191:184], PSPIC[0][183:176], PSPIC[0][175:168], PSPIC[0][167:160], PSPIC[0][159:152], PSPIC[0][151:144], PSPIC[0][143:136], PSPIC[0][135:128], PSPIC[0][127:120], PSPIC[0][119:112], PSPIC[0][111:104], PSPIC[0][103:96], PSPIC[0][95:88], PSPIC[0][87:80], PSPIC[0][79:72], PSPIC[0][71:64], PSPIC[0][63:56], PSPIC[0][55:48], PSPIC[0][47:40], PSPIC[0][39:32], PSPIC[0][31:24], PSPIC[0][23:16], PSPIC[0][15:8], PSPIC[0][7:0]};
assign PSPIC1 = { PSPIC[1][255:248], PSPIC[1][247:240], PSPIC[1][239:232], PSPIC[1][231:224], PSPIC[1][223:216], PSPIC[1][215:208], PSPIC[1][207:200], PSPIC[1][199:192], PSPIC[1][191:184], PSPIC[1][183:176], PSPIC[1][175:168], PSPIC[1][167:160], PSPIC[1][159:152], PSPIC[1][151:144], PSPIC[1][143:136], PSPIC[1][135:128], PSPIC[1][127:120], PSPIC[1][119:112], PSPIC[1][111:104], PSPIC[1][103:96], PSPIC[1][95:88], PSPIC[1][87:80], PSPIC[1][79:72], PSPIC[1][71:64], PSPIC[1][63:56], PSPIC[1][55:48], PSPIC[1][47:40], PSPIC[1][39:32], PSPIC[1][31:24], PSPIC[1][23:16], PSPIC[1][15:8], PSPIC[1][7:0]};
assign PSPIC2 = { PSPIC[2][255:248], PSPIC[2][247:240], PSPIC[2][239:232], PSPIC[2][231:224], PSPIC[2][223:216], PSPIC[2][215:208], PSPIC[2][207:200], PSPIC[2][199:192], PSPIC[2][191:184], PSPIC[2][183:176], PSPIC[2][175:168], PSPIC[2][167:160], PSPIC[2][159:152], PSPIC[2][151:144], PSPIC[2][143:136], PSPIC[2][135:128], PSPIC[2][127:120], PSPIC[2][119:112], PSPIC[2][111:104], PSPIC[2][103:96], PSPIC[2][95:88], PSPIC[2][87:80], PSPIC[2][79:72], PSPIC[2][71:64], PSPIC[2][63:56], PSPIC[2][55:48], PSPIC[2][47:40], PSPIC[2][39:32], PSPIC[2][31:24], PSPIC[2][23:16], PSPIC[2][15:8], PSPIC[2][7:0]};
assign PSPIC3 = { PSPIC[3][255:248], PSPIC[3][247:240], PSPIC[3][239:232], PSPIC[3][231:224], PSPIC[3][223:216], PSPIC[3][215:208], PSPIC[3][207:200], PSPIC[3][199:192], PSPIC[3][191:184], PSPIC[3][183:176], PSPIC[3][175:168], PSPIC[3][167:160], PSPIC[3][159:152], PSPIC[3][151:144], PSPIC[3][143:136], PSPIC[3][135:128], PSPIC[3][127:120], PSPIC[3][119:112], PSPIC[3][111:104], PSPIC[3][103:96], PSPIC[3][95:88], PSPIC[3][87:80], PSPIC[3][79:72], PSPIC[3][71:64], PSPIC[3][63:56], PSPIC[3][55:48], PSPIC[3][47:40], PSPIC[3][39:32], PSPIC[3][31:24], PSPIC[3][23:16], PSPIC[3][15:8], PSPIC[3][7:0]};
assign PSPIC4 = { PSPIC[4][255:248], PSPIC[4][247:240], PSPIC[4][239:232], PSPIC[4][231:224], PSPIC[4][223:216], PSPIC[4][215:208], PSPIC[4][207:200], PSPIC[4][199:192], PSPIC[4][191:184], PSPIC[4][183:176], PSPIC[4][175:168], PSPIC[4][167:160], PSPIC[4][159:152], PSPIC[4][151:144], PSPIC[4][143:136], PSPIC[4][135:128], PSPIC[4][127:120], PSPIC[4][119:112], PSPIC[4][111:104], PSPIC[4][103:96], PSPIC[4][95:88], PSPIC[4][87:80], PSPIC[4][79:72], PSPIC[4][71:64], PSPIC[4][63:56], PSPIC[4][55:48], PSPIC[4][47:40], PSPIC[4][39:32], PSPIC[4][31:24], PSPIC[4][23:16], PSPIC[4][15:8], PSPIC[4][7:0]};
assign PSPIC5 = { PSPIC[5][255:248], PSPIC[5][247:240], PSPIC[5][239:232], PSPIC[5][231:224], PSPIC[5][223:216], PSPIC[5][215:208], PSPIC[5][207:200], PSPIC[5][199:192], PSPIC[5][191:184], PSPIC[5][183:176], PSPIC[5][175:168], PSPIC[5][167:160], PSPIC[5][159:152], PSPIC[5][151:144], PSPIC[5][143:136], PSPIC[5][135:128], PSPIC[5][127:120], PSPIC[5][119:112], PSPIC[5][111:104], PSPIC[5][103:96], PSPIC[5][95:88], PSPIC[5][87:80], PSPIC[5][79:72], PSPIC[5][71:64], PSPIC[5][63:56], PSPIC[5][55:48], PSPIC[5][47:40], PSPIC[5][39:32], PSPIC[5][31:24], PSPIC[5][23:16], PSPIC[5][15:8], PSPIC[5][7:0]};
assign PSPIC6 = { PSPIC[6][255:248], PSPIC[6][247:240], PSPIC[6][239:232], PSPIC[6][231:224], PSPIC[6][223:216], PSPIC[6][215:208], PSPIC[6][207:200], PSPIC[6][199:192], PSPIC[6][191:184], PSPIC[6][183:176], PSPIC[6][175:168], PSPIC[6][167:160], PSPIC[6][159:152], PSPIC[6][151:144], PSPIC[6][143:136], PSPIC[6][135:128], PSPIC[6][127:120], PSPIC[6][119:112], PSPIC[6][111:104], PSPIC[6][103:96], PSPIC[6][95:88], PSPIC[6][87:80], PSPIC[6][79:72], PSPIC[6][71:64], PSPIC[6][63:56], PSPIC[6][55:48], PSPIC[6][47:40], PSPIC[6][39:32], PSPIC[6][31:24], PSPIC[6][23:16], PSPIC[6][15:8], PSPIC[6][7:0]};
assign PSPIC7 = { PSPIC[7][255:248], PSPIC[7][247:240], PSPIC[7][239:232], PSPIC[7][231:224], PSPIC[7][223:216], PSPIC[7][215:208], PSPIC[7][207:200], PSPIC[7][199:192], PSPIC[7][191:184], PSPIC[7][183:176], PSPIC[7][175:168], PSPIC[7][167:160], PSPIC[7][159:152], PSPIC[7][151:144], PSPIC[7][143:136], PSPIC[7][135:128], PSPIC[7][127:120], PSPIC[7][119:112], PSPIC[7][111:104], PSPIC[7][103:96], PSPIC[7][95:88], PSPIC[7][87:80], PSPIC[7][79:72], PSPIC[7][71:64], PSPIC[7][63:56], PSPIC[7][55:48], PSPIC[7][47:40], PSPIC[7][39:32], PSPIC[7][31:24], PSPIC[7][23:16], PSPIC[7][15:8], PSPIC[7][7:0]};
assign PSPIC8 = { PSPIC[8][255:248], PSPIC[8][247:240], PSPIC[8][239:232], PSPIC[8][231:224], PSPIC[8][223:216], PSPIC[8][215:208], PSPIC[8][207:200], PSPIC[8][199:192], PSPIC[8][191:184], PSPIC[8][183:176], PSPIC[8][175:168], PSPIC[8][167:160], PSPIC[8][159:152], PSPIC[8][151:144], PSPIC[8][143:136], PSPIC[8][135:128], PSPIC[8][127:120], PSPIC[8][119:112], PSPIC[8][111:104], PSPIC[8][103:96], PSPIC[8][95:88], PSPIC[8][87:80], PSPIC[8][79:72], PSPIC[8][71:64], PSPIC[8][63:56], PSPIC[8][55:48], PSPIC[8][47:40], PSPIC[8][39:32], PSPIC[8][31:24], PSPIC[8][23:16], PSPIC[8][15:8], PSPIC[8][7:0]};
assign PSPIC9 = { PSPIC[9][255:248], PSPIC[9][247:240], PSPIC[9][239:232], PSPIC[9][231:224], PSPIC[9][223:216], PSPIC[9][215:208], PSPIC[9][207:200], PSPIC[9][199:192], PSPIC[9][191:184], PSPIC[9][183:176], PSPIC[9][175:168], PSPIC[9][167:160], PSPIC[9][159:152], PSPIC[9][151:144], PSPIC[9][143:136], PSPIC[9][135:128], PSPIC[9][127:120], PSPIC[9][119:112], PSPIC[9][111:104], PSPIC[9][103:96], PSPIC[9][95:88], PSPIC[9][87:80], PSPIC[9][79:72], PSPIC[9][71:64], PSPIC[9][63:56], PSPIC[9][55:48], PSPIC[9][47:40], PSPIC[9][39:32], PSPIC[9][31:24], PSPIC[9][23:16], PSPIC[9][15:8], PSPIC[9][7:0]};
assign PSPIC10 = { PSPIC[10][255:248], PSPIC[10][247:240], PSPIC[10][239:232], PSPIC[10][231:224], PSPIC[10][223:216], PSPIC[10][215:208], PSPIC[10][207:200], PSPIC[10][199:192], PSPIC[10][191:184], PSPIC[10][183:176], PSPIC[10][175:168], PSPIC[10][167:160], PSPIC[10][159:152], PSPIC[10][151:144], PSPIC[10][143:136], PSPIC[10][135:128], PSPIC[10][127:120], PSPIC[10][119:112], PSPIC[10][111:104], PSPIC[10][103:96], PSPIC[10][95:88], PSPIC[10][87:80], PSPIC[10][79:72], PSPIC[10][71:64], PSPIC[10][63:56], PSPIC[10][55:48], PSPIC[10][47:40], PSPIC[10][39:32], PSPIC[10][31:24], PSPIC[10][23:16], PSPIC[10][15:8], PSPIC[10][7:0]};
assign PSPIC11 = { PSPIC[11][255:248], PSPIC[11][247:240], PSPIC[11][239:232], PSPIC[11][231:224], PSPIC[11][223:216], PSPIC[11][215:208], PSPIC[11][207:200], PSPIC[11][199:192], PSPIC[11][191:184], PSPIC[11][183:176], PSPIC[11][175:168], PSPIC[11][167:160], PSPIC[11][159:152], PSPIC[11][151:144], PSPIC[11][143:136], PSPIC[11][135:128], PSPIC[11][127:120], PSPIC[11][119:112], PSPIC[11][111:104], PSPIC[11][103:96], PSPIC[11][95:88], PSPIC[11][87:80], PSPIC[11][79:72], PSPIC[11][71:64], PSPIC[11][63:56], PSPIC[11][55:48], PSPIC[11][47:40], PSPIC[11][39:32], PSPIC[11][31:24], PSPIC[11][23:16], PSPIC[11][15:8], PSPIC[11][7:0]};
assign PSPIC12 = { PSPIC[12][255:248], PSPIC[12][247:240], PSPIC[12][239:232], PSPIC[12][231:224], PSPIC[12][223:216], PSPIC[12][215:208], PSPIC[12][207:200], PSPIC[12][199:192], PSPIC[12][191:184], PSPIC[12][183:176], PSPIC[12][175:168], PSPIC[12][167:160], PSPIC[12][159:152], PSPIC[12][151:144], PSPIC[12][143:136], PSPIC[12][135:128], PSPIC[12][127:120], PSPIC[12][119:112], PSPIC[12][111:104], PSPIC[12][103:96], PSPIC[12][95:88], PSPIC[12][87:80], PSPIC[12][79:72], PSPIC[12][71:64], PSPIC[12][63:56], PSPIC[12][55:48], PSPIC[12][47:40], PSPIC[12][39:32], PSPIC[12][31:24], PSPIC[12][23:16], PSPIC[12][15:8], PSPIC[12][7:0]};
assign PSPIC13 = { PSPIC[13][255:248], PSPIC[13][247:240], PSPIC[13][239:232], PSPIC[13][231:224], PSPIC[13][223:216], PSPIC[13][215:208], PSPIC[13][207:200], PSPIC[13][199:192], PSPIC[13][191:184], PSPIC[13][183:176], PSPIC[13][175:168], PSPIC[13][167:160], PSPIC[13][159:152], PSPIC[13][151:144], PSPIC[13][143:136], PSPIC[13][135:128], PSPIC[13][127:120], PSPIC[13][119:112], PSPIC[13][111:104], PSPIC[13][103:96], PSPIC[13][95:88], PSPIC[13][87:80], PSPIC[13][79:72], PSPIC[13][71:64], PSPIC[13][63:56], PSPIC[13][55:48], PSPIC[13][47:40], PSPIC[13][39:32], PSPIC[13][31:24], PSPIC[13][23:16], PSPIC[13][15:8], PSPIC[13][7:0]};
assign PSPIC14 = { PSPIC[14][255:248], PSPIC[14][247:240], PSPIC[14][239:232], PSPIC[14][231:224], PSPIC[14][223:216], PSPIC[14][215:208], PSPIC[14][207:200], PSPIC[14][199:192], PSPIC[14][191:184], PSPIC[14][183:176], PSPIC[14][175:168], PSPIC[14][167:160], PSPIC[14][159:152], PSPIC[14][151:144], PSPIC[14][143:136], PSPIC[14][135:128], PSPIC[14][127:120], PSPIC[14][119:112], PSPIC[14][111:104], PSPIC[14][103:96], PSPIC[14][95:88], PSPIC[14][87:80], PSPIC[14][79:72], PSPIC[14][71:64], PSPIC[14][63:56], PSPIC[14][55:48], PSPIC[14][47:40], PSPIC[14][39:32], PSPIC[14][31:24], PSPIC[14][23:16], PSPIC[14][15:8], PSPIC[14][7:0]};
assign PSPIC15 = { PSPIC[15][255:248], PSPIC[15][247:240], PSPIC[15][239:232], PSPIC[15][231:224], PSPIC[15][223:216], PSPIC[15][215:208], PSPIC[15][207:200], PSPIC[15][199:192], PSPIC[15][191:184], PSPIC[15][183:176], PSPIC[15][175:168], PSPIC[15][167:160], PSPIC[15][159:152], PSPIC[15][151:144], PSPIC[15][143:136], PSPIC[15][135:128], PSPIC[15][127:120], PSPIC[15][119:112], PSPIC[15][111:104], PSPIC[15][103:96], PSPIC[15][95:88], PSPIC[15][87:80], PSPIC[15][79:72], PSPIC[15][71:64], PSPIC[15][63:56], PSPIC[15][55:48], PSPIC[15][47:40], PSPIC[15][39:32], PSPIC[15][31:24], PSPIC[15][23:16], PSPIC[15][15:8], PSPIC[15][7:0]};
assign PSPIC16 = { PSPIC[16][255:248], PSPIC[16][247:240], PSPIC[16][239:232], PSPIC[16][231:224], PSPIC[16][223:216], PSPIC[16][215:208], PSPIC[16][207:200], PSPIC[16][199:192], PSPIC[16][191:184], PSPIC[16][183:176], PSPIC[16][175:168], PSPIC[16][167:160], PSPIC[16][159:152], PSPIC[16][151:144], PSPIC[16][143:136], PSPIC[16][135:128], PSPIC[16][127:120], PSPIC[16][119:112], PSPIC[16][111:104], PSPIC[16][103:96], PSPIC[16][95:88], PSPIC[16][87:80], PSPIC[16][79:72], PSPIC[16][71:64], PSPIC[16][63:56], PSPIC[16][55:48], PSPIC[16][47:40], PSPIC[16][39:32], PSPIC[16][31:24], PSPIC[16][23:16], PSPIC[16][15:8], PSPIC[16][7:0]};
assign PSPIC17 = { PSPIC[17][255:248], PSPIC[17][247:240], PSPIC[17][239:232], PSPIC[17][231:224], PSPIC[17][223:216], PSPIC[17][215:208], PSPIC[17][207:200], PSPIC[17][199:192], PSPIC[17][191:184], PSPIC[17][183:176], PSPIC[17][175:168], PSPIC[17][167:160], PSPIC[17][159:152], PSPIC[17][151:144], PSPIC[17][143:136], PSPIC[17][135:128], PSPIC[17][127:120], PSPIC[17][119:112], PSPIC[17][111:104], PSPIC[17][103:96], PSPIC[17][95:88], PSPIC[17][87:80], PSPIC[17][79:72], PSPIC[17][71:64], PSPIC[17][63:56], PSPIC[17][55:48], PSPIC[17][47:40], PSPIC[17][39:32], PSPIC[17][31:24], PSPIC[17][23:16], PSPIC[17][15:8], PSPIC[17][7:0]};
assign PSPIC18 = { PSPIC[18][255:248], PSPIC[18][247:240], PSPIC[18][239:232], PSPIC[18][231:224], PSPIC[18][223:216], PSPIC[18][215:208], PSPIC[18][207:200], PSPIC[18][199:192], PSPIC[18][191:184], PSPIC[18][183:176], PSPIC[18][175:168], PSPIC[18][167:160], PSPIC[18][159:152], PSPIC[18][151:144], PSPIC[18][143:136], PSPIC[18][135:128], PSPIC[18][127:120], PSPIC[18][119:112], PSPIC[18][111:104], PSPIC[18][103:96], PSPIC[18][95:88], PSPIC[18][87:80], PSPIC[18][79:72], PSPIC[18][71:64], PSPIC[18][63:56], PSPIC[18][55:48], PSPIC[18][47:40], PSPIC[18][39:32], PSPIC[18][31:24], PSPIC[18][23:16], PSPIC[18][15:8], PSPIC[18][7:0]};
assign PSPIC19 = { PSPIC[19][255:248], PSPIC[19][247:240], PSPIC[19][239:232], PSPIC[19][231:224], PSPIC[19][223:216], PSPIC[19][215:208], PSPIC[19][207:200], PSPIC[19][199:192], PSPIC[19][191:184], PSPIC[19][183:176], PSPIC[19][175:168], PSPIC[19][167:160], PSPIC[19][159:152], PSPIC[19][151:144], PSPIC[19][143:136], PSPIC[19][135:128], PSPIC[19][127:120], PSPIC[19][119:112], PSPIC[19][111:104], PSPIC[19][103:96], PSPIC[19][95:88], PSPIC[19][87:80], PSPIC[19][79:72], PSPIC[19][71:64], PSPIC[19][63:56], PSPIC[19][55:48], PSPIC[19][47:40], PSPIC[19][39:32], PSPIC[19][31:24], PSPIC[19][23:16], PSPIC[19][15:8], PSPIC[19][7:0]};
assign PSPIC20 = { PSPIC[20][255:248], PSPIC[20][247:240], PSPIC[20][239:232], PSPIC[20][231:224], PSPIC[20][223:216], PSPIC[20][215:208], PSPIC[20][207:200], PSPIC[20][199:192], PSPIC[20][191:184], PSPIC[20][183:176], PSPIC[20][175:168], PSPIC[20][167:160], PSPIC[20][159:152], PSPIC[20][151:144], PSPIC[20][143:136], PSPIC[20][135:128], PSPIC[20][127:120], PSPIC[20][119:112], PSPIC[20][111:104], PSPIC[20][103:96], PSPIC[20][95:88], PSPIC[20][87:80], PSPIC[20][79:72], PSPIC[20][71:64], PSPIC[20][63:56], PSPIC[20][55:48], PSPIC[20][47:40], PSPIC[20][39:32], PSPIC[20][31:24], PSPIC[20][23:16], PSPIC[20][15:8], PSPIC[20][7:0]};
assign PSPIC21 = { PSPIC[21][255:248], PSPIC[21][247:240], PSPIC[21][239:232], PSPIC[21][231:224], PSPIC[21][223:216], PSPIC[21][215:208], PSPIC[21][207:200], PSPIC[21][199:192], PSPIC[21][191:184], PSPIC[21][183:176], PSPIC[21][175:168], PSPIC[21][167:160], PSPIC[21][159:152], PSPIC[21][151:144], PSPIC[21][143:136], PSPIC[21][135:128], PSPIC[21][127:120], PSPIC[21][119:112], PSPIC[21][111:104], PSPIC[21][103:96], PSPIC[21][95:88], PSPIC[21][87:80], PSPIC[21][79:72], PSPIC[21][71:64], PSPIC[21][63:56], PSPIC[21][55:48], PSPIC[21][47:40], PSPIC[21][39:32], PSPIC[21][31:24], PSPIC[21][23:16], PSPIC[21][15:8], PSPIC[21][7:0]};
assign PSPIC22 = { PSPIC[22][255:248], PSPIC[22][247:240], PSPIC[22][239:232], PSPIC[22][231:224], PSPIC[22][223:216], PSPIC[22][215:208], PSPIC[22][207:200], PSPIC[22][199:192], PSPIC[22][191:184], PSPIC[22][183:176], PSPIC[22][175:168], PSPIC[22][167:160], PSPIC[22][159:152], PSPIC[22][151:144], PSPIC[22][143:136], PSPIC[22][135:128], PSPIC[22][127:120], PSPIC[22][119:112], PSPIC[22][111:104], PSPIC[22][103:96], PSPIC[22][95:88], PSPIC[22][87:80], PSPIC[22][79:72], PSPIC[22][71:64], PSPIC[22][63:56], PSPIC[22][55:48], PSPIC[22][47:40], PSPIC[22][39:32], PSPIC[22][31:24], PSPIC[22][23:16], PSPIC[22][15:8], PSPIC[22][7:0]};
assign PSPIC23 = { PSPIC[23][255:248], PSPIC[23][247:240], PSPIC[23][239:232], PSPIC[23][231:224], PSPIC[23][223:216], PSPIC[23][215:208], PSPIC[23][207:200], PSPIC[23][199:192], PSPIC[23][191:184], PSPIC[23][183:176], PSPIC[23][175:168], PSPIC[23][167:160], PSPIC[23][159:152], PSPIC[23][151:144], PSPIC[23][143:136], PSPIC[23][135:128], PSPIC[23][127:120], PSPIC[23][119:112], PSPIC[23][111:104], PSPIC[23][103:96], PSPIC[23][95:88], PSPIC[23][87:80], PSPIC[23][79:72], PSPIC[23][71:64], PSPIC[23][63:56], PSPIC[23][55:48], PSPIC[23][47:40], PSPIC[23][39:32], PSPIC[23][31:24], PSPIC[23][23:16], PSPIC[23][15:8], PSPIC[23][7:0]};
assign PSPIC24 = { PSPIC[24][255:248], PSPIC[24][247:240], PSPIC[24][239:232], PSPIC[24][231:224], PSPIC[24][223:216], PSPIC[24][215:208], PSPIC[24][207:200], PSPIC[24][199:192], PSPIC[24][191:184], PSPIC[24][183:176], PSPIC[24][175:168], PSPIC[24][167:160], PSPIC[24][159:152], PSPIC[24][151:144], PSPIC[24][143:136], PSPIC[24][135:128], PSPIC[24][127:120], PSPIC[24][119:112], PSPIC[24][111:104], PSPIC[24][103:96], PSPIC[24][95:88], PSPIC[24][87:80], PSPIC[24][79:72], PSPIC[24][71:64], PSPIC[24][63:56], PSPIC[24][55:48], PSPIC[24][47:40], PSPIC[24][39:32], PSPIC[24][31:24], PSPIC[24][23:16], PSPIC[24][15:8], PSPIC[24][7:0]};
assign PSPIC25 = { PSPIC[25][255:248], PSPIC[25][247:240], PSPIC[25][239:232], PSPIC[25][231:224], PSPIC[25][223:216], PSPIC[25][215:208], PSPIC[25][207:200], PSPIC[25][199:192], PSPIC[25][191:184], PSPIC[25][183:176], PSPIC[25][175:168], PSPIC[25][167:160], PSPIC[25][159:152], PSPIC[25][151:144], PSPIC[25][143:136], PSPIC[25][135:128], PSPIC[25][127:120], PSPIC[25][119:112], PSPIC[25][111:104], PSPIC[25][103:96], PSPIC[25][95:88], PSPIC[25][87:80], PSPIC[25][79:72], PSPIC[25][71:64], PSPIC[25][63:56], PSPIC[25][55:48], PSPIC[25][47:40], PSPIC[25][39:32], PSPIC[25][31:24], PSPIC[25][23:16], PSPIC[25][15:8], PSPIC[25][7:0]};
assign PSPIC26 = { PSPIC[26][255:248], PSPIC[26][247:240], PSPIC[26][239:232], PSPIC[26][231:224], PSPIC[26][223:216], PSPIC[26][215:208], PSPIC[26][207:200], PSPIC[26][199:192], PSPIC[26][191:184], PSPIC[26][183:176], PSPIC[26][175:168], PSPIC[26][167:160], PSPIC[26][159:152], PSPIC[26][151:144], PSPIC[26][143:136], PSPIC[26][135:128], PSPIC[26][127:120], PSPIC[26][119:112], PSPIC[26][111:104], PSPIC[26][103:96], PSPIC[26][95:88], PSPIC[26][87:80], PSPIC[26][79:72], PSPIC[26][71:64], PSPIC[26][63:56], PSPIC[26][55:48], PSPIC[26][47:40], PSPIC[26][39:32], PSPIC[26][31:24], PSPIC[26][23:16], PSPIC[26][15:8], PSPIC[26][7:0]};
assign PSPIC27 = { PSPIC[27][255:248], PSPIC[27][247:240], PSPIC[27][239:232], PSPIC[27][231:224], PSPIC[27][223:216], PSPIC[27][215:208], PSPIC[27][207:200], PSPIC[27][199:192], PSPIC[27][191:184], PSPIC[27][183:176], PSPIC[27][175:168], PSPIC[27][167:160], PSPIC[27][159:152], PSPIC[27][151:144], PSPIC[27][143:136], PSPIC[27][135:128], PSPIC[27][127:120], PSPIC[27][119:112], PSPIC[27][111:104], PSPIC[27][103:96], PSPIC[27][95:88], PSPIC[27][87:80], PSPIC[27][79:72], PSPIC[27][71:64], PSPIC[27][63:56], PSPIC[27][55:48], PSPIC[27][47:40], PSPIC[27][39:32], PSPIC[27][31:24], PSPIC[27][23:16], PSPIC[27][15:8], PSPIC[27][7:0]};
assign PSPIC28 = { PSPIC[28][255:248], PSPIC[28][247:240], PSPIC[28][239:232], PSPIC[28][231:224], PSPIC[28][223:216], PSPIC[28][215:208], PSPIC[28][207:200], PSPIC[28][199:192], PSPIC[28][191:184], PSPIC[28][183:176], PSPIC[28][175:168], PSPIC[28][167:160], PSPIC[28][159:152], PSPIC[28][151:144], PSPIC[28][143:136], PSPIC[28][135:128], PSPIC[28][127:120], PSPIC[28][119:112], PSPIC[28][111:104], PSPIC[28][103:96], PSPIC[28][95:88], PSPIC[28][87:80], PSPIC[28][79:72], PSPIC[28][71:64], PSPIC[28][63:56], PSPIC[28][55:48], PSPIC[28][47:40], PSPIC[28][39:32], PSPIC[28][31:24], PSPIC[28][23:16], PSPIC[28][15:8], PSPIC[28][7:0]};
assign PSPIC29 = { PSPIC[29][255:248], PSPIC[29][247:240], PSPIC[29][239:232], PSPIC[29][231:224], PSPIC[29][223:216], PSPIC[29][215:208], PSPIC[29][207:200], PSPIC[29][199:192], PSPIC[29][191:184], PSPIC[29][183:176], PSPIC[29][175:168], PSPIC[29][167:160], PSPIC[29][159:152], PSPIC[29][151:144], PSPIC[29][143:136], PSPIC[29][135:128], PSPIC[29][127:120], PSPIC[29][119:112], PSPIC[29][111:104], PSPIC[29][103:96], PSPIC[29][95:88], PSPIC[29][87:80], PSPIC[29][79:72], PSPIC[29][71:64], PSPIC[29][63:56], PSPIC[29][55:48], PSPIC[29][47:40], PSPIC[29][39:32], PSPIC[29][31:24], PSPIC[29][23:16], PSPIC[29][15:8], PSPIC[29][7:0]};
assign PSPIC30 = { PSPIC[30][255:248], PSPIC[30][247:240], PSPIC[30][239:232], PSPIC[30][231:224], PSPIC[30][223:216], PSPIC[30][215:208], PSPIC[30][207:200], PSPIC[30][199:192], PSPIC[30][191:184], PSPIC[30][183:176], PSPIC[30][175:168], PSPIC[30][167:160], PSPIC[30][159:152], PSPIC[30][151:144], PSPIC[30][143:136], PSPIC[30][135:128], PSPIC[30][127:120], PSPIC[30][119:112], PSPIC[30][111:104], PSPIC[30][103:96], PSPIC[30][95:88], PSPIC[30][87:80], PSPIC[30][79:72], PSPIC[30][71:64], PSPIC[30][63:56], PSPIC[30][55:48], PSPIC[30][47:40], PSPIC[30][39:32], PSPIC[30][31:24], PSPIC[30][23:16], PSPIC[30][15:8], PSPIC[30][7:0]};
assign PSPIC31 = { PSPIC[31][255:248], PSPIC[31][247:240], PSPIC[31][239:232], PSPIC[31][231:224], PSPIC[31][223:216], PSPIC[31][215:208], PSPIC[31][207:200], PSPIC[31][199:192], PSPIC[31][191:184], PSPIC[31][183:176], PSPIC[31][175:168], PSPIC[31][167:160], PSPIC[31][159:152], PSPIC[31][151:144], PSPIC[31][143:136], PSPIC[31][135:128], PSPIC[31][127:120], PSPIC[31][119:112], PSPIC[31][111:104], PSPIC[31][103:96], PSPIC[31][95:88], PSPIC[31][87:80], PSPIC[31][79:72], PSPIC[31][71:64], PSPIC[31][63:56], PSPIC[31][55:48], PSPIC[31][47:40], PSPIC[31][39:32], PSPIC[31][31:24], PSPIC[31][23:16], PSPIC[31][15:8], PSPIC[31][7:0]};




endmodule


